module mac5(a_t, a_f, a_ack, b_t, b_f, b_ack, out_t, out_f, out_ack, clk, reset);
input  clk, reset;
drwire csa_tree_add_14_36_groupi_n_0 ();
drwire csa_tree_add_14_36_groupi_n_1 ();
drwire csa_tree_add_14_36_groupi_n_10 ();
drwire csa_tree_add_14_36_groupi_n_100 ();
drwire csa_tree_add_14_36_groupi_n_1000 ();
drwire csa_tree_add_14_36_groupi_n_1001 ();
drwire csa_tree_add_14_36_groupi_n_1002 ();
drwire csa_tree_add_14_36_groupi_n_1003 ();
drwire csa_tree_add_14_36_groupi_n_1005 ();
drwire csa_tree_add_14_36_groupi_n_1006 ();
drwire csa_tree_add_14_36_groupi_n_1007 ();
drwire csa_tree_add_14_36_groupi_n_1008 ();
drwire csa_tree_add_14_36_groupi_n_1009 ();
drwire csa_tree_add_14_36_groupi_n_101 ();
drwire csa_tree_add_14_36_groupi_n_1010 ();
drwire csa_tree_add_14_36_groupi_n_1012 ();
drwire csa_tree_add_14_36_groupi_n_1013 ();
drwire csa_tree_add_14_36_groupi_n_1014 ();
drwire csa_tree_add_14_36_groupi_n_1015 ();
drwire csa_tree_add_14_36_groupi_n_1016 ();
drwire csa_tree_add_14_36_groupi_n_1017 ();
drwire csa_tree_add_14_36_groupi_n_1018 ();
drwire csa_tree_add_14_36_groupi_n_102 ();
drwire csa_tree_add_14_36_groupi_n_1020 ();
drwire csa_tree_add_14_36_groupi_n_1021 ();
drwire csa_tree_add_14_36_groupi_n_1022 ();
drwire csa_tree_add_14_36_groupi_n_1023 ();
drwire csa_tree_add_14_36_groupi_n_1024 ();
drwire csa_tree_add_14_36_groupi_n_1025 ();
drwire csa_tree_add_14_36_groupi_n_1026 ();
drwire csa_tree_add_14_36_groupi_n_1027 ();
drwire csa_tree_add_14_36_groupi_n_1028 ();
drwire csa_tree_add_14_36_groupi_n_1029 ();
drwire csa_tree_add_14_36_groupi_n_103 ();
drwire csa_tree_add_14_36_groupi_n_1030 ();
drwire csa_tree_add_14_36_groupi_n_1031 ();
drwire csa_tree_add_14_36_groupi_n_1032 ();
drwire csa_tree_add_14_36_groupi_n_1034 ();
drwire csa_tree_add_14_36_groupi_n_1036 ();
drwire csa_tree_add_14_36_groupi_n_1037 ();
drwire csa_tree_add_14_36_groupi_n_1038 ();
drwire csa_tree_add_14_36_groupi_n_1039 ();
drwire csa_tree_add_14_36_groupi_n_104 ();
drwire csa_tree_add_14_36_groupi_n_1040 ();
drwire csa_tree_add_14_36_groupi_n_1041 ();
drwire csa_tree_add_14_36_groupi_n_1042 ();
drwire csa_tree_add_14_36_groupi_n_1043 ();
drwire csa_tree_add_14_36_groupi_n_1044 ();
drwire csa_tree_add_14_36_groupi_n_1045 ();
drwire csa_tree_add_14_36_groupi_n_1046 ();
drwire csa_tree_add_14_36_groupi_n_1047 ();
drwire csa_tree_add_14_36_groupi_n_1048 ();
drwire csa_tree_add_14_36_groupi_n_1049 ();
drwire csa_tree_add_14_36_groupi_n_1050 ();
drwire csa_tree_add_14_36_groupi_n_1051 ();
drwire csa_tree_add_14_36_groupi_n_1052 ();
drwire csa_tree_add_14_36_groupi_n_1053 ();
drwire csa_tree_add_14_36_groupi_n_1054 ();
drwire csa_tree_add_14_36_groupi_n_1055 ();
drwire csa_tree_add_14_36_groupi_n_1056 ();
drwire csa_tree_add_14_36_groupi_n_1057 ();
drwire csa_tree_add_14_36_groupi_n_1058 ();
drwire csa_tree_add_14_36_groupi_n_1059 ();
drwire csa_tree_add_14_36_groupi_n_1060 ();
drwire csa_tree_add_14_36_groupi_n_1061 ();
drwire csa_tree_add_14_36_groupi_n_1062 ();
drwire csa_tree_add_14_36_groupi_n_1063 ();
drwire csa_tree_add_14_36_groupi_n_1064 ();
drwire csa_tree_add_14_36_groupi_n_1065 ();
drwire csa_tree_add_14_36_groupi_n_1066 ();
drwire csa_tree_add_14_36_groupi_n_1067 ();
drwire csa_tree_add_14_36_groupi_n_1068 ();
drwire csa_tree_add_14_36_groupi_n_1069 ();
drwire csa_tree_add_14_36_groupi_n_107 ();
drwire csa_tree_add_14_36_groupi_n_1070 ();
drwire csa_tree_add_14_36_groupi_n_1071 ();
drwire csa_tree_add_14_36_groupi_n_1072 ();
drwire csa_tree_add_14_36_groupi_n_1073 ();
drwire csa_tree_add_14_36_groupi_n_1074 ();
drwire csa_tree_add_14_36_groupi_n_1075 ();
drwire csa_tree_add_14_36_groupi_n_1076 ();
drwire csa_tree_add_14_36_groupi_n_1077 ();
drwire csa_tree_add_14_36_groupi_n_1078 ();
drwire csa_tree_add_14_36_groupi_n_1079 ();
drwire csa_tree_add_14_36_groupi_n_1080 ();
drwire csa_tree_add_14_36_groupi_n_1081 ();
drwire csa_tree_add_14_36_groupi_n_1082 ();
drwire csa_tree_add_14_36_groupi_n_1083 ();
drwire csa_tree_add_14_36_groupi_n_1084 ();
drwire csa_tree_add_14_36_groupi_n_1085 ();
drwire csa_tree_add_14_36_groupi_n_1086 ();
drwire csa_tree_add_14_36_groupi_n_1087 ();
drwire csa_tree_add_14_36_groupi_n_1088 ();
drwire csa_tree_add_14_36_groupi_n_1089 ();
drwire csa_tree_add_14_36_groupi_n_109 ();
drwire csa_tree_add_14_36_groupi_n_1090 ();
drwire csa_tree_add_14_36_groupi_n_1092 ();
drwire csa_tree_add_14_36_groupi_n_1093 ();
drwire csa_tree_add_14_36_groupi_n_1094 ();
drwire csa_tree_add_14_36_groupi_n_1095 ();
drwire csa_tree_add_14_36_groupi_n_1096 ();
drwire csa_tree_add_14_36_groupi_n_1097 ();
drwire csa_tree_add_14_36_groupi_n_1098 ();
drwire csa_tree_add_14_36_groupi_n_1099 ();
drwire csa_tree_add_14_36_groupi_n_11 ();
drwire csa_tree_add_14_36_groupi_n_110 ();
drwire csa_tree_add_14_36_groupi_n_1100 ();
drwire csa_tree_add_14_36_groupi_n_1101 ();
drwire csa_tree_add_14_36_groupi_n_1102 ();
drwire csa_tree_add_14_36_groupi_n_1104 ();
drwire csa_tree_add_14_36_groupi_n_1105 ();
drwire csa_tree_add_14_36_groupi_n_1106 ();
drwire csa_tree_add_14_36_groupi_n_1107 ();
drwire csa_tree_add_14_36_groupi_n_1108 ();
drwire csa_tree_add_14_36_groupi_n_1109 ();
drwire csa_tree_add_14_36_groupi_n_1110 ();
drwire csa_tree_add_14_36_groupi_n_1111 ();
drwire csa_tree_add_14_36_groupi_n_1112 ();
drwire csa_tree_add_14_36_groupi_n_1113 ();
drwire csa_tree_add_14_36_groupi_n_1114 ();
drwire csa_tree_add_14_36_groupi_n_1115 ();
drwire csa_tree_add_14_36_groupi_n_1116 ();
drwire csa_tree_add_14_36_groupi_n_1118 ();
drwire csa_tree_add_14_36_groupi_n_1119 ();
drwire csa_tree_add_14_36_groupi_n_112 ();
drwire csa_tree_add_14_36_groupi_n_1120 ();
drwire csa_tree_add_14_36_groupi_n_1121 ();
drwire csa_tree_add_14_36_groupi_n_1122 ();
drwire csa_tree_add_14_36_groupi_n_1123 ();
drwire csa_tree_add_14_36_groupi_n_1125 ();
drwire csa_tree_add_14_36_groupi_n_1126 ();
drwire csa_tree_add_14_36_groupi_n_1127 ();
drwire csa_tree_add_14_36_groupi_n_1128 ();
drwire csa_tree_add_14_36_groupi_n_113 ();
drwire csa_tree_add_14_36_groupi_n_1130 ();
drwire csa_tree_add_14_36_groupi_n_1132 ();
drwire csa_tree_add_14_36_groupi_n_1133 ();
drwire csa_tree_add_14_36_groupi_n_1135 ();
drwire csa_tree_add_14_36_groupi_n_1136 ();
drwire csa_tree_add_14_36_groupi_n_1137 ();
drwire csa_tree_add_14_36_groupi_n_1138 ();
drwire csa_tree_add_14_36_groupi_n_1139 ();
drwire csa_tree_add_14_36_groupi_n_114 ();
drwire csa_tree_add_14_36_groupi_n_1140 ();
drwire csa_tree_add_14_36_groupi_n_1141 ();
drwire csa_tree_add_14_36_groupi_n_1142 ();
drwire csa_tree_add_14_36_groupi_n_1144 ();
drwire csa_tree_add_14_36_groupi_n_1146 ();
drwire csa_tree_add_14_36_groupi_n_1147 ();
drwire csa_tree_add_14_36_groupi_n_1148 ();
drwire csa_tree_add_14_36_groupi_n_1149 ();
drwire csa_tree_add_14_36_groupi_n_115 ();
drwire csa_tree_add_14_36_groupi_n_1151 ();
drwire csa_tree_add_14_36_groupi_n_1152 ();
drwire csa_tree_add_14_36_groupi_n_1153 ();
drwire csa_tree_add_14_36_groupi_n_1154 ();
drwire csa_tree_add_14_36_groupi_n_1155 ();
drwire csa_tree_add_14_36_groupi_n_116 ();
drwire csa_tree_add_14_36_groupi_n_1160 ();
drwire csa_tree_add_14_36_groupi_n_1162 ();
drwire csa_tree_add_14_36_groupi_n_1163 ();
drwire csa_tree_add_14_36_groupi_n_1164 ();
drwire csa_tree_add_14_36_groupi_n_1165 ();
drwire csa_tree_add_14_36_groupi_n_1166 ();
drwire csa_tree_add_14_36_groupi_n_1167 ();
drwire csa_tree_add_14_36_groupi_n_1168 ();
drwire csa_tree_add_14_36_groupi_n_1169 ();
drwire csa_tree_add_14_36_groupi_n_117 ();
drwire csa_tree_add_14_36_groupi_n_1170 ();
drwire csa_tree_add_14_36_groupi_n_1171 ();
drwire csa_tree_add_14_36_groupi_n_1172 ();
drwire csa_tree_add_14_36_groupi_n_1174 ();
drwire csa_tree_add_14_36_groupi_n_1175 ();
drwire csa_tree_add_14_36_groupi_n_1177 ();
drwire csa_tree_add_14_36_groupi_n_1178 ();
drwire csa_tree_add_14_36_groupi_n_1179 ();
drwire csa_tree_add_14_36_groupi_n_118 ();
drwire csa_tree_add_14_36_groupi_n_1180 ();
drwire csa_tree_add_14_36_groupi_n_1181 ();
drwire csa_tree_add_14_36_groupi_n_1184 ();
drwire csa_tree_add_14_36_groupi_n_1185 ();
drwire csa_tree_add_14_36_groupi_n_1186 ();
drwire csa_tree_add_14_36_groupi_n_1187 ();
drwire csa_tree_add_14_36_groupi_n_1188 ();
drwire csa_tree_add_14_36_groupi_n_1189 ();
drwire csa_tree_add_14_36_groupi_n_119 ();
drwire csa_tree_add_14_36_groupi_n_1190 ();
drwire csa_tree_add_14_36_groupi_n_1191 ();
drwire csa_tree_add_14_36_groupi_n_1192 ();
drwire csa_tree_add_14_36_groupi_n_1193 ();
drwire csa_tree_add_14_36_groupi_n_1195 ();
drwire csa_tree_add_14_36_groupi_n_1196 ();
drwire csa_tree_add_14_36_groupi_n_1197 ();
drwire csa_tree_add_14_36_groupi_n_1198 ();
drwire csa_tree_add_14_36_groupi_n_1199 ();
drwire csa_tree_add_14_36_groupi_n_120 ();
drwire csa_tree_add_14_36_groupi_n_1200 ();
drwire csa_tree_add_14_36_groupi_n_1201 ();
drwire csa_tree_add_14_36_groupi_n_1202 ();
drwire csa_tree_add_14_36_groupi_n_1203 ();
drwire csa_tree_add_14_36_groupi_n_1204 ();
drwire csa_tree_add_14_36_groupi_n_1205 ();
drwire csa_tree_add_14_36_groupi_n_1206 ();
drwire csa_tree_add_14_36_groupi_n_1209 ();
drwire csa_tree_add_14_36_groupi_n_121 ();
drwire csa_tree_add_14_36_groupi_n_1210 ();
drwire csa_tree_add_14_36_groupi_n_1211 ();
drwire csa_tree_add_14_36_groupi_n_1212 ();
drwire csa_tree_add_14_36_groupi_n_1214 ();
drwire csa_tree_add_14_36_groupi_n_1215 ();
drwire csa_tree_add_14_36_groupi_n_1216 ();
drwire csa_tree_add_14_36_groupi_n_1217 ();
drwire csa_tree_add_14_36_groupi_n_1219 ();
drwire csa_tree_add_14_36_groupi_n_122 ();
drwire csa_tree_add_14_36_groupi_n_1221 ();
drwire csa_tree_add_14_36_groupi_n_1222 ();
drwire csa_tree_add_14_36_groupi_n_1223 ();
drwire csa_tree_add_14_36_groupi_n_1224 ();
drwire csa_tree_add_14_36_groupi_n_1225 ();
drwire csa_tree_add_14_36_groupi_n_1226 ();
drwire csa_tree_add_14_36_groupi_n_1227 ();
drwire csa_tree_add_14_36_groupi_n_1228 ();
drwire csa_tree_add_14_36_groupi_n_1229 ();
drwire csa_tree_add_14_36_groupi_n_123 ();
drwire csa_tree_add_14_36_groupi_n_1230 ();
drwire csa_tree_add_14_36_groupi_n_1231 ();
drwire csa_tree_add_14_36_groupi_n_1232 ();
drwire csa_tree_add_14_36_groupi_n_1234 ();
drwire csa_tree_add_14_36_groupi_n_1235 ();
drwire csa_tree_add_14_36_groupi_n_1236 ();
drwire csa_tree_add_14_36_groupi_n_1237 ();
drwire csa_tree_add_14_36_groupi_n_1238 ();
drwire csa_tree_add_14_36_groupi_n_1239 ();
drwire csa_tree_add_14_36_groupi_n_124 ();
drwire csa_tree_add_14_36_groupi_n_1241 ();
drwire csa_tree_add_14_36_groupi_n_1242 ();
drwire csa_tree_add_14_36_groupi_n_1243 ();
drwire csa_tree_add_14_36_groupi_n_1245 ();
drwire csa_tree_add_14_36_groupi_n_1246 ();
drwire csa_tree_add_14_36_groupi_n_1247 ();
drwire csa_tree_add_14_36_groupi_n_1248 ();
drwire csa_tree_add_14_36_groupi_n_1249 ();
drwire csa_tree_add_14_36_groupi_n_125 ();
drwire csa_tree_add_14_36_groupi_n_1250 ();
drwire csa_tree_add_14_36_groupi_n_1251 ();
drwire csa_tree_add_14_36_groupi_n_1252 ();
drwire csa_tree_add_14_36_groupi_n_1253 ();
drwire csa_tree_add_14_36_groupi_n_1254 ();
drwire csa_tree_add_14_36_groupi_n_1255 ();
drwire csa_tree_add_14_36_groupi_n_1256 ();
drwire csa_tree_add_14_36_groupi_n_1257 ();
drwire csa_tree_add_14_36_groupi_n_1258 ();
drwire csa_tree_add_14_36_groupi_n_1259 ();
drwire csa_tree_add_14_36_groupi_n_1260 ();
drwire csa_tree_add_14_36_groupi_n_1261 ();
drwire csa_tree_add_14_36_groupi_n_1262 ();
drwire csa_tree_add_14_36_groupi_n_1263 ();
drwire csa_tree_add_14_36_groupi_n_1264 ();
drwire csa_tree_add_14_36_groupi_n_1265 ();
drwire csa_tree_add_14_36_groupi_n_1266 ();
drwire csa_tree_add_14_36_groupi_n_1267 ();
drwire csa_tree_add_14_36_groupi_n_1269 ();
drwire csa_tree_add_14_36_groupi_n_127 ();
drwire csa_tree_add_14_36_groupi_n_1270 ();
drwire csa_tree_add_14_36_groupi_n_1272 ();
drwire csa_tree_add_14_36_groupi_n_1273 ();
drwire csa_tree_add_14_36_groupi_n_1274 ();
drwire csa_tree_add_14_36_groupi_n_1275 ();
drwire csa_tree_add_14_36_groupi_n_1276 ();
drwire csa_tree_add_14_36_groupi_n_1278 ();
drwire csa_tree_add_14_36_groupi_n_1279 ();
drwire csa_tree_add_14_36_groupi_n_128 ();
drwire csa_tree_add_14_36_groupi_n_1280 ();
drwire csa_tree_add_14_36_groupi_n_1281 ();
drwire csa_tree_add_14_36_groupi_n_1282 ();
drwire csa_tree_add_14_36_groupi_n_1283 ();
drwire csa_tree_add_14_36_groupi_n_1284 ();
drwire csa_tree_add_14_36_groupi_n_1285 ();
drwire csa_tree_add_14_36_groupi_n_1286 ();
drwire csa_tree_add_14_36_groupi_n_1287 ();
drwire csa_tree_add_14_36_groupi_n_1288 ();
drwire csa_tree_add_14_36_groupi_n_1289 ();
drwire csa_tree_add_14_36_groupi_n_129 ();
drwire csa_tree_add_14_36_groupi_n_1290 ();
drwire csa_tree_add_14_36_groupi_n_1291 ();
drwire csa_tree_add_14_36_groupi_n_1292 ();
drwire csa_tree_add_14_36_groupi_n_1293 ();
drwire csa_tree_add_14_36_groupi_n_1294 ();
drwire csa_tree_add_14_36_groupi_n_1295 ();
drwire csa_tree_add_14_36_groupi_n_1296 ();
drwire csa_tree_add_14_36_groupi_n_1299 ();
drwire csa_tree_add_14_36_groupi_n_13 ();
drwire csa_tree_add_14_36_groupi_n_130 ();
drwire csa_tree_add_14_36_groupi_n_1300 ();
drwire csa_tree_add_14_36_groupi_n_1301 ();
drwire csa_tree_add_14_36_groupi_n_1302 ();
drwire csa_tree_add_14_36_groupi_n_1303 ();
drwire csa_tree_add_14_36_groupi_n_1304 ();
drwire csa_tree_add_14_36_groupi_n_1305 ();
drwire csa_tree_add_14_36_groupi_n_1308 ();
drwire csa_tree_add_14_36_groupi_n_1309 ();
drwire csa_tree_add_14_36_groupi_n_1311 ();
drwire csa_tree_add_14_36_groupi_n_1312 ();
drwire csa_tree_add_14_36_groupi_n_1313 ();
drwire csa_tree_add_14_36_groupi_n_1314 ();
drwire csa_tree_add_14_36_groupi_n_1315 ();
drwire csa_tree_add_14_36_groupi_n_1316 ();
drwire csa_tree_add_14_36_groupi_n_1317 ();
drwire csa_tree_add_14_36_groupi_n_1318 ();
drwire csa_tree_add_14_36_groupi_n_1319 ();
drwire csa_tree_add_14_36_groupi_n_1320 ();
drwire csa_tree_add_14_36_groupi_n_1321 ();
drwire csa_tree_add_14_36_groupi_n_1322 ();
drwire csa_tree_add_14_36_groupi_n_1325 ();
drwire csa_tree_add_14_36_groupi_n_1326 ();
drwire csa_tree_add_14_36_groupi_n_1327 ();
drwire csa_tree_add_14_36_groupi_n_1329 ();
drwire csa_tree_add_14_36_groupi_n_1330 ();
drwire csa_tree_add_14_36_groupi_n_1331 ();
drwire csa_tree_add_14_36_groupi_n_1332 ();
drwire csa_tree_add_14_36_groupi_n_1333 ();
drwire csa_tree_add_14_36_groupi_n_1334 ();
drwire csa_tree_add_14_36_groupi_n_1335 ();
drwire csa_tree_add_14_36_groupi_n_1336 ();
drwire csa_tree_add_14_36_groupi_n_1337 ();
drwire csa_tree_add_14_36_groupi_n_1338 ();
drwire csa_tree_add_14_36_groupi_n_1339 ();
drwire csa_tree_add_14_36_groupi_n_134 ();
drwire csa_tree_add_14_36_groupi_n_1340 ();
drwire csa_tree_add_14_36_groupi_n_1341 ();
drwire csa_tree_add_14_36_groupi_n_1342 ();
drwire csa_tree_add_14_36_groupi_n_1343 ();
drwire csa_tree_add_14_36_groupi_n_1344 ();
drwire csa_tree_add_14_36_groupi_n_1345 ();
drwire csa_tree_add_14_36_groupi_n_1346 ();
drwire csa_tree_add_14_36_groupi_n_1347 ();
drwire csa_tree_add_14_36_groupi_n_1349 ();
drwire csa_tree_add_14_36_groupi_n_135 ();
drwire csa_tree_add_14_36_groupi_n_1350 ();
drwire csa_tree_add_14_36_groupi_n_1351 ();
drwire csa_tree_add_14_36_groupi_n_1352 ();
drwire csa_tree_add_14_36_groupi_n_1353 ();
drwire csa_tree_add_14_36_groupi_n_1354 ();
drwire csa_tree_add_14_36_groupi_n_1355 ();
drwire csa_tree_add_14_36_groupi_n_1356 ();
drwire csa_tree_add_14_36_groupi_n_1357 ();
drwire csa_tree_add_14_36_groupi_n_1358 ();
drwire csa_tree_add_14_36_groupi_n_1359 ();
drwire csa_tree_add_14_36_groupi_n_136 ();
drwire csa_tree_add_14_36_groupi_n_1361 ();
drwire csa_tree_add_14_36_groupi_n_1362 ();
drwire csa_tree_add_14_36_groupi_n_1363 ();
drwire csa_tree_add_14_36_groupi_n_1364 ();
drwire csa_tree_add_14_36_groupi_n_1365 ();
drwire csa_tree_add_14_36_groupi_n_1366 ();
drwire csa_tree_add_14_36_groupi_n_1367 ();
drwire csa_tree_add_14_36_groupi_n_1368 ();
drwire csa_tree_add_14_36_groupi_n_1369 ();
drwire csa_tree_add_14_36_groupi_n_137 ();
drwire csa_tree_add_14_36_groupi_n_1370 ();
drwire csa_tree_add_14_36_groupi_n_1371 ();
drwire csa_tree_add_14_36_groupi_n_1372 ();
drwire csa_tree_add_14_36_groupi_n_1373 ();
drwire csa_tree_add_14_36_groupi_n_1374 ();
drwire csa_tree_add_14_36_groupi_n_1375 ();
drwire csa_tree_add_14_36_groupi_n_1376 ();
drwire csa_tree_add_14_36_groupi_n_1377 ();
drwire csa_tree_add_14_36_groupi_n_1378 ();
drwire csa_tree_add_14_36_groupi_n_1379 ();
drwire csa_tree_add_14_36_groupi_n_138 ();
drwire csa_tree_add_14_36_groupi_n_1380 ();
drwire csa_tree_add_14_36_groupi_n_1381 ();
drwire csa_tree_add_14_36_groupi_n_1382 ();
drwire csa_tree_add_14_36_groupi_n_1383 ();
drwire csa_tree_add_14_36_groupi_n_1384 ();
drwire csa_tree_add_14_36_groupi_n_1385 ();
drwire csa_tree_add_14_36_groupi_n_1386 ();
drwire csa_tree_add_14_36_groupi_n_1387 ();
drwire csa_tree_add_14_36_groupi_n_1388 ();
drwire csa_tree_add_14_36_groupi_n_1389 ();
drwire csa_tree_add_14_36_groupi_n_139 ();
drwire csa_tree_add_14_36_groupi_n_1390 ();
drwire csa_tree_add_14_36_groupi_n_1391 ();
drwire csa_tree_add_14_36_groupi_n_1392 ();
drwire csa_tree_add_14_36_groupi_n_1393 ();
drwire csa_tree_add_14_36_groupi_n_1395 ();
drwire csa_tree_add_14_36_groupi_n_1396 ();
drwire csa_tree_add_14_36_groupi_n_1397 ();
drwire csa_tree_add_14_36_groupi_n_1398 ();
drwire csa_tree_add_14_36_groupi_n_1399 ();
drwire csa_tree_add_14_36_groupi_n_14 ();
drwire csa_tree_add_14_36_groupi_n_140 ();
drwire csa_tree_add_14_36_groupi_n_1400 ();
drwire csa_tree_add_14_36_groupi_n_1401 ();
drwire csa_tree_add_14_36_groupi_n_1402 ();
drwire csa_tree_add_14_36_groupi_n_1403 ();
drwire csa_tree_add_14_36_groupi_n_1405 ();
drwire csa_tree_add_14_36_groupi_n_1406 ();
drwire csa_tree_add_14_36_groupi_n_1407 ();
drwire csa_tree_add_14_36_groupi_n_1408 ();
drwire csa_tree_add_14_36_groupi_n_141 ();
drwire csa_tree_add_14_36_groupi_n_1411 ();
drwire csa_tree_add_14_36_groupi_n_1412 ();
drwire csa_tree_add_14_36_groupi_n_1413 ();
drwire csa_tree_add_14_36_groupi_n_1414 ();
drwire csa_tree_add_14_36_groupi_n_1415 ();
drwire csa_tree_add_14_36_groupi_n_1416 ();
drwire csa_tree_add_14_36_groupi_n_1417 ();
drwire csa_tree_add_14_36_groupi_n_1418 ();
drwire csa_tree_add_14_36_groupi_n_1419 ();
drwire csa_tree_add_14_36_groupi_n_142 ();
drwire csa_tree_add_14_36_groupi_n_1420 ();
drwire csa_tree_add_14_36_groupi_n_1421 ();
drwire csa_tree_add_14_36_groupi_n_1422 ();
drwire csa_tree_add_14_36_groupi_n_1423 ();
drwire csa_tree_add_14_36_groupi_n_1424 ();
drwire csa_tree_add_14_36_groupi_n_1425 ();
drwire csa_tree_add_14_36_groupi_n_1427 ();
drwire csa_tree_add_14_36_groupi_n_1428 ();
drwire csa_tree_add_14_36_groupi_n_1429 ();
drwire csa_tree_add_14_36_groupi_n_1430 ();
drwire csa_tree_add_14_36_groupi_n_1431 ();
drwire csa_tree_add_14_36_groupi_n_1432 ();
drwire csa_tree_add_14_36_groupi_n_1433 ();
drwire csa_tree_add_14_36_groupi_n_1434 ();
drwire csa_tree_add_14_36_groupi_n_1435 ();
drwire csa_tree_add_14_36_groupi_n_1436 ();
drwire csa_tree_add_14_36_groupi_n_1437 ();
drwire csa_tree_add_14_36_groupi_n_1438 ();
drwire csa_tree_add_14_36_groupi_n_1439 ();
drwire csa_tree_add_14_36_groupi_n_144 ();
drwire csa_tree_add_14_36_groupi_n_1440 ();
drwire csa_tree_add_14_36_groupi_n_1441 ();
drwire csa_tree_add_14_36_groupi_n_1442 ();
drwire csa_tree_add_14_36_groupi_n_1444 ();
drwire csa_tree_add_14_36_groupi_n_1445 ();
drwire csa_tree_add_14_36_groupi_n_1446 ();
drwire csa_tree_add_14_36_groupi_n_1447 ();
drwire csa_tree_add_14_36_groupi_n_1448 ();
drwire csa_tree_add_14_36_groupi_n_1449 ();
drwire csa_tree_add_14_36_groupi_n_1450 ();
drwire csa_tree_add_14_36_groupi_n_1451 ();
drwire csa_tree_add_14_36_groupi_n_1452 ();
drwire csa_tree_add_14_36_groupi_n_1453 ();
drwire csa_tree_add_14_36_groupi_n_1455 ();
drwire csa_tree_add_14_36_groupi_n_1456 ();
drwire csa_tree_add_14_36_groupi_n_1457 ();
drwire csa_tree_add_14_36_groupi_n_1458 ();
drwire csa_tree_add_14_36_groupi_n_1459 ();
drwire csa_tree_add_14_36_groupi_n_146 ();
drwire csa_tree_add_14_36_groupi_n_1460 ();
drwire csa_tree_add_14_36_groupi_n_1461 ();
drwire csa_tree_add_14_36_groupi_n_1462 ();
drwire csa_tree_add_14_36_groupi_n_1463 ();
drwire csa_tree_add_14_36_groupi_n_1464 ();
drwire csa_tree_add_14_36_groupi_n_1465 ();
drwire csa_tree_add_14_36_groupi_n_1466 ();
drwire csa_tree_add_14_36_groupi_n_1467 ();
drwire csa_tree_add_14_36_groupi_n_1468 ();
drwire csa_tree_add_14_36_groupi_n_147 ();
drwire csa_tree_add_14_36_groupi_n_1470 ();
drwire csa_tree_add_14_36_groupi_n_1471 ();
drwire csa_tree_add_14_36_groupi_n_1472 ();
drwire csa_tree_add_14_36_groupi_n_1473 ();
drwire csa_tree_add_14_36_groupi_n_1474 ();
drwire csa_tree_add_14_36_groupi_n_1475 ();
drwire csa_tree_add_14_36_groupi_n_1476 ();
drwire csa_tree_add_14_36_groupi_n_1477 ();
drwire csa_tree_add_14_36_groupi_n_1478 ();
drwire csa_tree_add_14_36_groupi_n_1479 ();
drwire csa_tree_add_14_36_groupi_n_148 ();
drwire csa_tree_add_14_36_groupi_n_1480 ();
drwire csa_tree_add_14_36_groupi_n_1481 ();
drwire csa_tree_add_14_36_groupi_n_1482 ();
drwire csa_tree_add_14_36_groupi_n_1483 ();
drwire csa_tree_add_14_36_groupi_n_1484 ();
drwire csa_tree_add_14_36_groupi_n_1485 ();
drwire csa_tree_add_14_36_groupi_n_1486 ();
drwire csa_tree_add_14_36_groupi_n_1487 ();
drwire csa_tree_add_14_36_groupi_n_1488 ();
drwire csa_tree_add_14_36_groupi_n_1489 ();
drwire csa_tree_add_14_36_groupi_n_1490 ();
drwire csa_tree_add_14_36_groupi_n_1491 ();
drwire csa_tree_add_14_36_groupi_n_1492 ();
drwire csa_tree_add_14_36_groupi_n_1493 ();
drwire csa_tree_add_14_36_groupi_n_1494 ();
drwire csa_tree_add_14_36_groupi_n_1495 ();
drwire csa_tree_add_14_36_groupi_n_1496 ();
drwire csa_tree_add_14_36_groupi_n_1497 ();
drwire csa_tree_add_14_36_groupi_n_1498 ();
drwire csa_tree_add_14_36_groupi_n_1499 ();
drwire csa_tree_add_14_36_groupi_n_15 ();
drwire csa_tree_add_14_36_groupi_n_150 ();
drwire csa_tree_add_14_36_groupi_n_1500 ();
drwire csa_tree_add_14_36_groupi_n_1501 ();
drwire csa_tree_add_14_36_groupi_n_1502 ();
drwire csa_tree_add_14_36_groupi_n_1503 ();
drwire csa_tree_add_14_36_groupi_n_1504 ();
drwire csa_tree_add_14_36_groupi_n_1505 ();
drwire csa_tree_add_14_36_groupi_n_1506 ();
drwire csa_tree_add_14_36_groupi_n_1507 ();
drwire csa_tree_add_14_36_groupi_n_1508 ();
drwire csa_tree_add_14_36_groupi_n_1509 ();
drwire csa_tree_add_14_36_groupi_n_151 ();
drwire csa_tree_add_14_36_groupi_n_1510 ();
drwire csa_tree_add_14_36_groupi_n_1512 ();
drwire csa_tree_add_14_36_groupi_n_1513 ();
drwire csa_tree_add_14_36_groupi_n_1514 ();
drwire csa_tree_add_14_36_groupi_n_1516 ();
drwire csa_tree_add_14_36_groupi_n_1517 ();
drwire csa_tree_add_14_36_groupi_n_1518 ();
drwire csa_tree_add_14_36_groupi_n_1519 ();
drwire csa_tree_add_14_36_groupi_n_152 ();
drwire csa_tree_add_14_36_groupi_n_1520 ();
drwire csa_tree_add_14_36_groupi_n_1521 ();
drwire csa_tree_add_14_36_groupi_n_1522 ();
drwire csa_tree_add_14_36_groupi_n_1523 ();
drwire csa_tree_add_14_36_groupi_n_1524 ();
drwire csa_tree_add_14_36_groupi_n_1525 ();
drwire csa_tree_add_14_36_groupi_n_1526 ();
drwire csa_tree_add_14_36_groupi_n_1527 ();
drwire csa_tree_add_14_36_groupi_n_1528 ();
drwire csa_tree_add_14_36_groupi_n_1529 ();
drwire csa_tree_add_14_36_groupi_n_153 ();
drwire csa_tree_add_14_36_groupi_n_1530 ();
drwire csa_tree_add_14_36_groupi_n_1531 ();
drwire csa_tree_add_14_36_groupi_n_1532 ();
drwire csa_tree_add_14_36_groupi_n_1533 ();
drwire csa_tree_add_14_36_groupi_n_1534 ();
drwire csa_tree_add_14_36_groupi_n_1535 ();
drwire csa_tree_add_14_36_groupi_n_1536 ();
drwire csa_tree_add_14_36_groupi_n_1537 ();
drwire csa_tree_add_14_36_groupi_n_1538 ();
drwire csa_tree_add_14_36_groupi_n_1539 ();
drwire csa_tree_add_14_36_groupi_n_154 ();
drwire csa_tree_add_14_36_groupi_n_1540 ();
drwire csa_tree_add_14_36_groupi_n_1541 ();
drwire csa_tree_add_14_36_groupi_n_1542 ();
drwire csa_tree_add_14_36_groupi_n_1543 ();
drwire csa_tree_add_14_36_groupi_n_1547 ();
drwire csa_tree_add_14_36_groupi_n_1548 ();
drwire csa_tree_add_14_36_groupi_n_1549 ();
drwire csa_tree_add_14_36_groupi_n_155 ();
drwire csa_tree_add_14_36_groupi_n_1550 ();
drwire csa_tree_add_14_36_groupi_n_1551 ();
drwire csa_tree_add_14_36_groupi_n_1552 ();
drwire csa_tree_add_14_36_groupi_n_1553 ();
drwire csa_tree_add_14_36_groupi_n_1554 ();
drwire csa_tree_add_14_36_groupi_n_1555 ();
drwire csa_tree_add_14_36_groupi_n_1556 ();
drwire csa_tree_add_14_36_groupi_n_1557 ();
drwire csa_tree_add_14_36_groupi_n_1558 ();
drwire csa_tree_add_14_36_groupi_n_1559 ();
drwire csa_tree_add_14_36_groupi_n_156 ();
drwire csa_tree_add_14_36_groupi_n_1560 ();
drwire csa_tree_add_14_36_groupi_n_1561 ();
drwire csa_tree_add_14_36_groupi_n_1562 ();
drwire csa_tree_add_14_36_groupi_n_1563 ();
drwire csa_tree_add_14_36_groupi_n_1564 ();
drwire csa_tree_add_14_36_groupi_n_1565 ();
drwire csa_tree_add_14_36_groupi_n_1566 ();
drwire csa_tree_add_14_36_groupi_n_1567 ();
drwire csa_tree_add_14_36_groupi_n_1568 ();
drwire csa_tree_add_14_36_groupi_n_1569 ();
drwire csa_tree_add_14_36_groupi_n_157 ();
drwire csa_tree_add_14_36_groupi_n_1571 ();
drwire csa_tree_add_14_36_groupi_n_1572 ();
drwire csa_tree_add_14_36_groupi_n_1573 ();
drwire csa_tree_add_14_36_groupi_n_1574 ();
drwire csa_tree_add_14_36_groupi_n_1575 ();
drwire csa_tree_add_14_36_groupi_n_1577 ();
drwire csa_tree_add_14_36_groupi_n_1578 ();
drwire csa_tree_add_14_36_groupi_n_1579 ();
drwire csa_tree_add_14_36_groupi_n_158 ();
drwire csa_tree_add_14_36_groupi_n_1580 ();
drwire csa_tree_add_14_36_groupi_n_1581 ();
drwire csa_tree_add_14_36_groupi_n_1582 ();
drwire csa_tree_add_14_36_groupi_n_1583 ();
drwire csa_tree_add_14_36_groupi_n_1584 ();
drwire csa_tree_add_14_36_groupi_n_1585 ();
drwire csa_tree_add_14_36_groupi_n_1586 ();
drwire csa_tree_add_14_36_groupi_n_1587 ();
drwire csa_tree_add_14_36_groupi_n_1588 ();
drwire csa_tree_add_14_36_groupi_n_1589 ();
drwire csa_tree_add_14_36_groupi_n_159 ();
drwire csa_tree_add_14_36_groupi_n_1590 ();
drwire csa_tree_add_14_36_groupi_n_1591 ();
drwire csa_tree_add_14_36_groupi_n_1594 ();
drwire csa_tree_add_14_36_groupi_n_1595 ();
drwire csa_tree_add_14_36_groupi_n_1596 ();
drwire csa_tree_add_14_36_groupi_n_1597 ();
drwire csa_tree_add_14_36_groupi_n_1598 ();
drwire csa_tree_add_14_36_groupi_n_1599 ();
drwire csa_tree_add_14_36_groupi_n_16 ();
drwire csa_tree_add_14_36_groupi_n_160 ();
drwire csa_tree_add_14_36_groupi_n_1600 ();
drwire csa_tree_add_14_36_groupi_n_1601 ();
drwire csa_tree_add_14_36_groupi_n_1602 ();
drwire csa_tree_add_14_36_groupi_n_1604 ();
drwire csa_tree_add_14_36_groupi_n_1605 ();
drwire csa_tree_add_14_36_groupi_n_1607 ();
drwire csa_tree_add_14_36_groupi_n_1608 ();
drwire csa_tree_add_14_36_groupi_n_1609 ();
drwire csa_tree_add_14_36_groupi_n_161 ();
drwire csa_tree_add_14_36_groupi_n_1610 ();
drwire csa_tree_add_14_36_groupi_n_1611 ();
drwire csa_tree_add_14_36_groupi_n_1612 ();
drwire csa_tree_add_14_36_groupi_n_1613 ();
drwire csa_tree_add_14_36_groupi_n_1614 ();
drwire csa_tree_add_14_36_groupi_n_1615 ();
drwire csa_tree_add_14_36_groupi_n_1616 ();
drwire csa_tree_add_14_36_groupi_n_1617 ();
drwire csa_tree_add_14_36_groupi_n_1618 ();
drwire csa_tree_add_14_36_groupi_n_1619 ();
drwire csa_tree_add_14_36_groupi_n_162 ();
drwire csa_tree_add_14_36_groupi_n_1620 ();
drwire csa_tree_add_14_36_groupi_n_1621 ();
drwire csa_tree_add_14_36_groupi_n_1622 ();
drwire csa_tree_add_14_36_groupi_n_1623 ();
drwire csa_tree_add_14_36_groupi_n_1624 ();
drwire csa_tree_add_14_36_groupi_n_1625 ();
drwire csa_tree_add_14_36_groupi_n_1627 ();
drwire csa_tree_add_14_36_groupi_n_1629 ();
drwire csa_tree_add_14_36_groupi_n_163 ();
drwire csa_tree_add_14_36_groupi_n_1630 ();
drwire csa_tree_add_14_36_groupi_n_1631 ();
drwire csa_tree_add_14_36_groupi_n_1633 ();
drwire csa_tree_add_14_36_groupi_n_1634 ();
drwire csa_tree_add_14_36_groupi_n_1635 ();
drwire csa_tree_add_14_36_groupi_n_1636 ();
drwire csa_tree_add_14_36_groupi_n_1637 ();
drwire csa_tree_add_14_36_groupi_n_1639 ();
drwire csa_tree_add_14_36_groupi_n_164 ();
drwire csa_tree_add_14_36_groupi_n_1640 ();
drwire csa_tree_add_14_36_groupi_n_1642 ();
drwire csa_tree_add_14_36_groupi_n_1643 ();
drwire csa_tree_add_14_36_groupi_n_1644 ();
drwire csa_tree_add_14_36_groupi_n_1645 ();
drwire csa_tree_add_14_36_groupi_n_1646 ();
drwire csa_tree_add_14_36_groupi_n_1647 ();
drwire csa_tree_add_14_36_groupi_n_1648 ();
drwire csa_tree_add_14_36_groupi_n_1649 ();
drwire csa_tree_add_14_36_groupi_n_165 ();
drwire csa_tree_add_14_36_groupi_n_1650 ();
drwire csa_tree_add_14_36_groupi_n_1651 ();
drwire csa_tree_add_14_36_groupi_n_1652 ();
drwire csa_tree_add_14_36_groupi_n_1653 ();
drwire csa_tree_add_14_36_groupi_n_1654 ();
drwire csa_tree_add_14_36_groupi_n_1655 ();
drwire csa_tree_add_14_36_groupi_n_1656 ();
drwire csa_tree_add_14_36_groupi_n_1657 ();
drwire csa_tree_add_14_36_groupi_n_166 ();
drwire csa_tree_add_14_36_groupi_n_1661 ();
drwire csa_tree_add_14_36_groupi_n_1662 ();
drwire csa_tree_add_14_36_groupi_n_1663 ();
drwire csa_tree_add_14_36_groupi_n_1664 ();
drwire csa_tree_add_14_36_groupi_n_1666 ();
drwire csa_tree_add_14_36_groupi_n_1667 ();
drwire csa_tree_add_14_36_groupi_n_1668 ();
drwire csa_tree_add_14_36_groupi_n_1669 ();
drwire csa_tree_add_14_36_groupi_n_167 ();
drwire csa_tree_add_14_36_groupi_n_1670 ();
drwire csa_tree_add_14_36_groupi_n_1671 ();
drwire csa_tree_add_14_36_groupi_n_1672 ();
drwire csa_tree_add_14_36_groupi_n_1673 ();
drwire csa_tree_add_14_36_groupi_n_1674 ();
drwire csa_tree_add_14_36_groupi_n_1676 ();
drwire csa_tree_add_14_36_groupi_n_1677 ();
drwire csa_tree_add_14_36_groupi_n_1678 ();
drwire csa_tree_add_14_36_groupi_n_1679 ();
drwire csa_tree_add_14_36_groupi_n_168 ();
drwire csa_tree_add_14_36_groupi_n_1680 ();
drwire csa_tree_add_14_36_groupi_n_1681 ();
drwire csa_tree_add_14_36_groupi_n_1682 ();
drwire csa_tree_add_14_36_groupi_n_1683 ();
drwire csa_tree_add_14_36_groupi_n_1684 ();
drwire csa_tree_add_14_36_groupi_n_1685 ();
drwire csa_tree_add_14_36_groupi_n_1686 ();
drwire csa_tree_add_14_36_groupi_n_1687 ();
drwire csa_tree_add_14_36_groupi_n_1688 ();
drwire csa_tree_add_14_36_groupi_n_169 ();
drwire csa_tree_add_14_36_groupi_n_1690 ();
drwire csa_tree_add_14_36_groupi_n_1691 ();
drwire csa_tree_add_14_36_groupi_n_1693 ();
drwire csa_tree_add_14_36_groupi_n_1694 ();
drwire csa_tree_add_14_36_groupi_n_1695 ();
drwire csa_tree_add_14_36_groupi_n_1696 ();
drwire csa_tree_add_14_36_groupi_n_1697 ();
drwire csa_tree_add_14_36_groupi_n_1698 ();
drwire csa_tree_add_14_36_groupi_n_1699 ();
drwire csa_tree_add_14_36_groupi_n_17 ();
drwire csa_tree_add_14_36_groupi_n_170 ();
drwire csa_tree_add_14_36_groupi_n_1700 ();
drwire csa_tree_add_14_36_groupi_n_1701 ();
drwire csa_tree_add_14_36_groupi_n_1702 ();
drwire csa_tree_add_14_36_groupi_n_1703 ();
drwire csa_tree_add_14_36_groupi_n_1704 ();
drwire csa_tree_add_14_36_groupi_n_1705 ();
drwire csa_tree_add_14_36_groupi_n_1706 ();
drwire csa_tree_add_14_36_groupi_n_1707 ();
drwire csa_tree_add_14_36_groupi_n_1708 ();
drwire csa_tree_add_14_36_groupi_n_1709 ();
drwire csa_tree_add_14_36_groupi_n_171 ();
drwire csa_tree_add_14_36_groupi_n_1710 ();
drwire csa_tree_add_14_36_groupi_n_1711 ();
drwire csa_tree_add_14_36_groupi_n_1712 ();
drwire csa_tree_add_14_36_groupi_n_1713 ();
drwire csa_tree_add_14_36_groupi_n_1714 ();
drwire csa_tree_add_14_36_groupi_n_1715 ();
drwire csa_tree_add_14_36_groupi_n_1716 ();
drwire csa_tree_add_14_36_groupi_n_1717 ();
drwire csa_tree_add_14_36_groupi_n_1718 ();
drwire csa_tree_add_14_36_groupi_n_1719 ();
drwire csa_tree_add_14_36_groupi_n_172 ();
drwire csa_tree_add_14_36_groupi_n_1720 ();
drwire csa_tree_add_14_36_groupi_n_1721 ();
drwire csa_tree_add_14_36_groupi_n_1722 ();
drwire csa_tree_add_14_36_groupi_n_1723 ();
drwire csa_tree_add_14_36_groupi_n_1724 ();
drwire csa_tree_add_14_36_groupi_n_1725 ();
drwire csa_tree_add_14_36_groupi_n_1726 ();
drwire csa_tree_add_14_36_groupi_n_1727 ();
drwire csa_tree_add_14_36_groupi_n_1728 ();
drwire csa_tree_add_14_36_groupi_n_1729 ();
drwire csa_tree_add_14_36_groupi_n_173 ();
drwire csa_tree_add_14_36_groupi_n_1730 ();
drwire csa_tree_add_14_36_groupi_n_1731 ();
drwire csa_tree_add_14_36_groupi_n_1733 ();
drwire csa_tree_add_14_36_groupi_n_1734 ();
drwire csa_tree_add_14_36_groupi_n_1735 ();
drwire csa_tree_add_14_36_groupi_n_1737 ();
drwire csa_tree_add_14_36_groupi_n_1738 ();
drwire csa_tree_add_14_36_groupi_n_174 ();
drwire csa_tree_add_14_36_groupi_n_1740 ();
drwire csa_tree_add_14_36_groupi_n_1741 ();
drwire csa_tree_add_14_36_groupi_n_1742 ();
drwire csa_tree_add_14_36_groupi_n_1743 ();
drwire csa_tree_add_14_36_groupi_n_1744 ();
drwire csa_tree_add_14_36_groupi_n_1746 ();
drwire csa_tree_add_14_36_groupi_n_1747 ();
drwire csa_tree_add_14_36_groupi_n_1748 ();
drwire csa_tree_add_14_36_groupi_n_1749 ();
drwire csa_tree_add_14_36_groupi_n_175 ();
drwire csa_tree_add_14_36_groupi_n_1751 ();
drwire csa_tree_add_14_36_groupi_n_1753 ();
drwire csa_tree_add_14_36_groupi_n_1754 ();
drwire csa_tree_add_14_36_groupi_n_1756 ();
drwire csa_tree_add_14_36_groupi_n_1757 ();
drwire csa_tree_add_14_36_groupi_n_1758 ();
drwire csa_tree_add_14_36_groupi_n_176 ();
drwire csa_tree_add_14_36_groupi_n_1760 ();
drwire csa_tree_add_14_36_groupi_n_1761 ();
drwire csa_tree_add_14_36_groupi_n_1762 ();
drwire csa_tree_add_14_36_groupi_n_1763 ();
drwire csa_tree_add_14_36_groupi_n_1764 ();
drwire csa_tree_add_14_36_groupi_n_1765 ();
drwire csa_tree_add_14_36_groupi_n_1766 ();
drwire csa_tree_add_14_36_groupi_n_1767 ();
drwire csa_tree_add_14_36_groupi_n_1768 ();
drwire csa_tree_add_14_36_groupi_n_1769 ();
drwire csa_tree_add_14_36_groupi_n_177 ();
drwire csa_tree_add_14_36_groupi_n_1770 ();
drwire csa_tree_add_14_36_groupi_n_1771 ();
drwire csa_tree_add_14_36_groupi_n_1772 ();
drwire csa_tree_add_14_36_groupi_n_1773 ();
drwire csa_tree_add_14_36_groupi_n_1774 ();
drwire csa_tree_add_14_36_groupi_n_1775 ();
drwire csa_tree_add_14_36_groupi_n_1776 ();
drwire csa_tree_add_14_36_groupi_n_1777 ();
drwire csa_tree_add_14_36_groupi_n_1778 ();
drwire csa_tree_add_14_36_groupi_n_1779 ();
drwire csa_tree_add_14_36_groupi_n_178 ();
drwire csa_tree_add_14_36_groupi_n_1780 ();
drwire csa_tree_add_14_36_groupi_n_1781 ();
drwire csa_tree_add_14_36_groupi_n_1782 ();
drwire csa_tree_add_14_36_groupi_n_1785 ();
drwire csa_tree_add_14_36_groupi_n_1786 ();
drwire csa_tree_add_14_36_groupi_n_1787 ();
drwire csa_tree_add_14_36_groupi_n_1788 ();
drwire csa_tree_add_14_36_groupi_n_1789 ();
drwire csa_tree_add_14_36_groupi_n_179 ();
drwire csa_tree_add_14_36_groupi_n_1790 ();
drwire csa_tree_add_14_36_groupi_n_1791 ();
drwire csa_tree_add_14_36_groupi_n_1792 ();
drwire csa_tree_add_14_36_groupi_n_1793 ();
drwire csa_tree_add_14_36_groupi_n_1794 ();
drwire csa_tree_add_14_36_groupi_n_1795 ();
drwire csa_tree_add_14_36_groupi_n_1796 ();
drwire csa_tree_add_14_36_groupi_n_1797 ();
drwire csa_tree_add_14_36_groupi_n_1798 ();
drwire csa_tree_add_14_36_groupi_n_1799 ();
drwire csa_tree_add_14_36_groupi_n_18 ();
drwire csa_tree_add_14_36_groupi_n_180 ();
drwire csa_tree_add_14_36_groupi_n_1800 ();
drwire csa_tree_add_14_36_groupi_n_1801 ();
drwire csa_tree_add_14_36_groupi_n_1802 ();
drwire csa_tree_add_14_36_groupi_n_1803 ();
drwire csa_tree_add_14_36_groupi_n_1804 ();
drwire csa_tree_add_14_36_groupi_n_1805 ();
drwire csa_tree_add_14_36_groupi_n_1806 ();
drwire csa_tree_add_14_36_groupi_n_1807 ();
drwire csa_tree_add_14_36_groupi_n_1808 ();
drwire csa_tree_add_14_36_groupi_n_1809 ();
drwire csa_tree_add_14_36_groupi_n_181 ();
drwire csa_tree_add_14_36_groupi_n_1810 ();
drwire csa_tree_add_14_36_groupi_n_1811 ();
drwire csa_tree_add_14_36_groupi_n_1812 ();
drwire csa_tree_add_14_36_groupi_n_1813 ();
drwire csa_tree_add_14_36_groupi_n_1814 ();
drwire csa_tree_add_14_36_groupi_n_1815 ();
drwire csa_tree_add_14_36_groupi_n_1816 ();
drwire csa_tree_add_14_36_groupi_n_1817 ();
drwire csa_tree_add_14_36_groupi_n_1818 ();
drwire csa_tree_add_14_36_groupi_n_1819 ();
drwire csa_tree_add_14_36_groupi_n_182 ();
drwire csa_tree_add_14_36_groupi_n_1820 ();
drwire csa_tree_add_14_36_groupi_n_1821 ();
drwire csa_tree_add_14_36_groupi_n_1822 ();
drwire csa_tree_add_14_36_groupi_n_1823 ();
drwire csa_tree_add_14_36_groupi_n_1824 ();
drwire csa_tree_add_14_36_groupi_n_1825 ();
drwire csa_tree_add_14_36_groupi_n_1826 ();
drwire csa_tree_add_14_36_groupi_n_1827 ();
drwire csa_tree_add_14_36_groupi_n_1828 ();
drwire csa_tree_add_14_36_groupi_n_1829 ();
drwire csa_tree_add_14_36_groupi_n_183 ();
drwire csa_tree_add_14_36_groupi_n_1830 ();
drwire csa_tree_add_14_36_groupi_n_1831 ();
drwire csa_tree_add_14_36_groupi_n_1832 ();
drwire csa_tree_add_14_36_groupi_n_1833 ();
drwire csa_tree_add_14_36_groupi_n_1834 ();
drwire csa_tree_add_14_36_groupi_n_1835 ();
drwire csa_tree_add_14_36_groupi_n_1836 ();
drwire csa_tree_add_14_36_groupi_n_1837 ();
drwire csa_tree_add_14_36_groupi_n_1838 ();
drwire csa_tree_add_14_36_groupi_n_1839 ();
drwire csa_tree_add_14_36_groupi_n_184 ();
drwire csa_tree_add_14_36_groupi_n_1840 ();
drwire csa_tree_add_14_36_groupi_n_1841 ();
drwire csa_tree_add_14_36_groupi_n_1842 ();
drwire csa_tree_add_14_36_groupi_n_1843 ();
drwire csa_tree_add_14_36_groupi_n_1844 ();
drwire csa_tree_add_14_36_groupi_n_1845 ();
drwire csa_tree_add_14_36_groupi_n_1846 ();
drwire csa_tree_add_14_36_groupi_n_1847 ();
drwire csa_tree_add_14_36_groupi_n_1848 ();
drwire csa_tree_add_14_36_groupi_n_1849 ();
drwire csa_tree_add_14_36_groupi_n_185 ();
drwire csa_tree_add_14_36_groupi_n_1850 ();
drwire csa_tree_add_14_36_groupi_n_1851 ();
drwire csa_tree_add_14_36_groupi_n_1853 ();
drwire csa_tree_add_14_36_groupi_n_1854 ();
drwire csa_tree_add_14_36_groupi_n_1855 ();
drwire csa_tree_add_14_36_groupi_n_1856 ();
drwire csa_tree_add_14_36_groupi_n_1857 ();
drwire csa_tree_add_14_36_groupi_n_1858 ();
drwire csa_tree_add_14_36_groupi_n_1859 ();
drwire csa_tree_add_14_36_groupi_n_186 ();
drwire csa_tree_add_14_36_groupi_n_1860 ();
drwire csa_tree_add_14_36_groupi_n_1861 ();
drwire csa_tree_add_14_36_groupi_n_1862 ();
drwire csa_tree_add_14_36_groupi_n_1863 ();
drwire csa_tree_add_14_36_groupi_n_1864 ();
drwire csa_tree_add_14_36_groupi_n_1865 ();
drwire csa_tree_add_14_36_groupi_n_1866 ();
drwire csa_tree_add_14_36_groupi_n_1867 ();
drwire csa_tree_add_14_36_groupi_n_1868 ();
drwire csa_tree_add_14_36_groupi_n_1869 ();
drwire csa_tree_add_14_36_groupi_n_187 ();
drwire csa_tree_add_14_36_groupi_n_1870 ();
drwire csa_tree_add_14_36_groupi_n_1871 ();
drwire csa_tree_add_14_36_groupi_n_1873 ();
drwire csa_tree_add_14_36_groupi_n_1875 ();
drwire csa_tree_add_14_36_groupi_n_1876 ();
drwire csa_tree_add_14_36_groupi_n_1877 ();
drwire csa_tree_add_14_36_groupi_n_1878 ();
drwire csa_tree_add_14_36_groupi_n_1879 ();
drwire csa_tree_add_14_36_groupi_n_188 ();
drwire csa_tree_add_14_36_groupi_n_1880 ();
drwire csa_tree_add_14_36_groupi_n_1881 ();
drwire csa_tree_add_14_36_groupi_n_1882 ();
drwire csa_tree_add_14_36_groupi_n_1883 ();
drwire csa_tree_add_14_36_groupi_n_1884 ();
drwire csa_tree_add_14_36_groupi_n_1885 ();
drwire csa_tree_add_14_36_groupi_n_1886 ();
drwire csa_tree_add_14_36_groupi_n_1887 ();
drwire csa_tree_add_14_36_groupi_n_1888 ();
drwire csa_tree_add_14_36_groupi_n_1889 ();
drwire csa_tree_add_14_36_groupi_n_189 ();
drwire csa_tree_add_14_36_groupi_n_1890 ();
drwire csa_tree_add_14_36_groupi_n_1891 ();
drwire csa_tree_add_14_36_groupi_n_1892 ();
drwire csa_tree_add_14_36_groupi_n_1894 ();
drwire csa_tree_add_14_36_groupi_n_1895 ();
drwire csa_tree_add_14_36_groupi_n_1896 ();
drwire csa_tree_add_14_36_groupi_n_1897 ();
drwire csa_tree_add_14_36_groupi_n_1898 ();
drwire csa_tree_add_14_36_groupi_n_1899 ();
drwire csa_tree_add_14_36_groupi_n_19 ();
drwire csa_tree_add_14_36_groupi_n_190 ();
drwire csa_tree_add_14_36_groupi_n_1900 ();
drwire csa_tree_add_14_36_groupi_n_1901 ();
drwire csa_tree_add_14_36_groupi_n_1902 ();
drwire csa_tree_add_14_36_groupi_n_1903 ();
drwire csa_tree_add_14_36_groupi_n_1904 ();
drwire csa_tree_add_14_36_groupi_n_1905 ();
drwire csa_tree_add_14_36_groupi_n_1906 ();
drwire csa_tree_add_14_36_groupi_n_1907 ();
drwire csa_tree_add_14_36_groupi_n_1908 ();
drwire csa_tree_add_14_36_groupi_n_1909 ();
drwire csa_tree_add_14_36_groupi_n_191 ();
drwire csa_tree_add_14_36_groupi_n_1910 ();
drwire csa_tree_add_14_36_groupi_n_1911 ();
drwire csa_tree_add_14_36_groupi_n_1912 ();
drwire csa_tree_add_14_36_groupi_n_1913 ();
drwire csa_tree_add_14_36_groupi_n_1914 ();
drwire csa_tree_add_14_36_groupi_n_1915 ();
drwire csa_tree_add_14_36_groupi_n_1916 ();
drwire csa_tree_add_14_36_groupi_n_1917 ();
drwire csa_tree_add_14_36_groupi_n_1918 ();
drwire csa_tree_add_14_36_groupi_n_1919 ();
drwire csa_tree_add_14_36_groupi_n_192 ();
drwire csa_tree_add_14_36_groupi_n_1920 ();
drwire csa_tree_add_14_36_groupi_n_1921 ();
drwire csa_tree_add_14_36_groupi_n_1922 ();
drwire csa_tree_add_14_36_groupi_n_1923 ();
drwire csa_tree_add_14_36_groupi_n_1924 ();
drwire csa_tree_add_14_36_groupi_n_1925 ();
drwire csa_tree_add_14_36_groupi_n_1926 ();
drwire csa_tree_add_14_36_groupi_n_1927 ();
drwire csa_tree_add_14_36_groupi_n_1928 ();
drwire csa_tree_add_14_36_groupi_n_1929 ();
drwire csa_tree_add_14_36_groupi_n_193 ();
drwire csa_tree_add_14_36_groupi_n_1930 ();
drwire csa_tree_add_14_36_groupi_n_1931 ();
drwire csa_tree_add_14_36_groupi_n_1932 ();
drwire csa_tree_add_14_36_groupi_n_1933 ();
drwire csa_tree_add_14_36_groupi_n_1934 ();
drwire csa_tree_add_14_36_groupi_n_1935 ();
drwire csa_tree_add_14_36_groupi_n_1936 ();
drwire csa_tree_add_14_36_groupi_n_1937 ();
drwire csa_tree_add_14_36_groupi_n_1938 ();
drwire csa_tree_add_14_36_groupi_n_1939 ();
drwire csa_tree_add_14_36_groupi_n_194 ();
drwire csa_tree_add_14_36_groupi_n_1940 ();
drwire csa_tree_add_14_36_groupi_n_1941 ();
drwire csa_tree_add_14_36_groupi_n_1942 ();
drwire csa_tree_add_14_36_groupi_n_1943 ();
drwire csa_tree_add_14_36_groupi_n_1944 ();
drwire csa_tree_add_14_36_groupi_n_1945 ();
drwire csa_tree_add_14_36_groupi_n_1946 ();
drwire csa_tree_add_14_36_groupi_n_1947 ();
drwire csa_tree_add_14_36_groupi_n_1948 ();
drwire csa_tree_add_14_36_groupi_n_1949 ();
drwire csa_tree_add_14_36_groupi_n_195 ();
drwire csa_tree_add_14_36_groupi_n_1950 ();
drwire csa_tree_add_14_36_groupi_n_1951 ();
drwire csa_tree_add_14_36_groupi_n_1952 ();
drwire csa_tree_add_14_36_groupi_n_1953 ();
drwire csa_tree_add_14_36_groupi_n_1954 ();
drwire csa_tree_add_14_36_groupi_n_1955 ();
drwire csa_tree_add_14_36_groupi_n_1956 ();
drwire csa_tree_add_14_36_groupi_n_1957 ();
drwire csa_tree_add_14_36_groupi_n_1958 ();
drwire csa_tree_add_14_36_groupi_n_1959 ();
drwire csa_tree_add_14_36_groupi_n_196 ();
drwire csa_tree_add_14_36_groupi_n_1960 ();
drwire csa_tree_add_14_36_groupi_n_1961 ();
drwire csa_tree_add_14_36_groupi_n_1962 ();
drwire csa_tree_add_14_36_groupi_n_1963 ();
drwire csa_tree_add_14_36_groupi_n_1964 ();
drwire csa_tree_add_14_36_groupi_n_1965 ();
drwire csa_tree_add_14_36_groupi_n_1966 ();
drwire csa_tree_add_14_36_groupi_n_1967 ();
drwire csa_tree_add_14_36_groupi_n_1968 ();
drwire csa_tree_add_14_36_groupi_n_1969 ();
drwire csa_tree_add_14_36_groupi_n_197 ();
drwire csa_tree_add_14_36_groupi_n_1970 ();
drwire csa_tree_add_14_36_groupi_n_1971 ();
drwire csa_tree_add_14_36_groupi_n_1972 ();
drwire csa_tree_add_14_36_groupi_n_1973 ();
drwire csa_tree_add_14_36_groupi_n_1974 ();
drwire csa_tree_add_14_36_groupi_n_1975 ();
drwire csa_tree_add_14_36_groupi_n_1976 ();
drwire csa_tree_add_14_36_groupi_n_1977 ();
drwire csa_tree_add_14_36_groupi_n_1978 ();
drwire csa_tree_add_14_36_groupi_n_1979 ();
drwire csa_tree_add_14_36_groupi_n_198 ();
drwire csa_tree_add_14_36_groupi_n_1980 ();
drwire csa_tree_add_14_36_groupi_n_1981 ();
drwire csa_tree_add_14_36_groupi_n_1982 ();
drwire csa_tree_add_14_36_groupi_n_1983 ();
drwire csa_tree_add_14_36_groupi_n_1984 ();
drwire csa_tree_add_14_36_groupi_n_1985 ();
drwire csa_tree_add_14_36_groupi_n_1986 ();
drwire csa_tree_add_14_36_groupi_n_1987 ();
drwire csa_tree_add_14_36_groupi_n_1988 ();
drwire csa_tree_add_14_36_groupi_n_1989 ();
drwire csa_tree_add_14_36_groupi_n_199 ();
drwire csa_tree_add_14_36_groupi_n_1990 ();
drwire csa_tree_add_14_36_groupi_n_1991 ();
drwire csa_tree_add_14_36_groupi_n_1992 ();
drwire csa_tree_add_14_36_groupi_n_1993 ();
drwire csa_tree_add_14_36_groupi_n_1994 ();
drwire csa_tree_add_14_36_groupi_n_1995 ();
drwire csa_tree_add_14_36_groupi_n_1996 ();
drwire csa_tree_add_14_36_groupi_n_1997 ();
drwire csa_tree_add_14_36_groupi_n_1998 ();
drwire csa_tree_add_14_36_groupi_n_1999 ();
drwire csa_tree_add_14_36_groupi_n_2 ();
drwire csa_tree_add_14_36_groupi_n_20 ();
drwire csa_tree_add_14_36_groupi_n_200 ();
drwire csa_tree_add_14_36_groupi_n_2000 ();
drwire csa_tree_add_14_36_groupi_n_2001 ();
drwire csa_tree_add_14_36_groupi_n_2002 ();
drwire csa_tree_add_14_36_groupi_n_2003 ();
drwire csa_tree_add_14_36_groupi_n_2004 ();
drwire csa_tree_add_14_36_groupi_n_2005 ();
drwire csa_tree_add_14_36_groupi_n_2006 ();
drwire csa_tree_add_14_36_groupi_n_2007 ();
drwire csa_tree_add_14_36_groupi_n_2008 ();
drwire csa_tree_add_14_36_groupi_n_2009 ();
drwire csa_tree_add_14_36_groupi_n_201 ();
drwire csa_tree_add_14_36_groupi_n_2010 ();
drwire csa_tree_add_14_36_groupi_n_2011 ();
drwire csa_tree_add_14_36_groupi_n_2012 ();
drwire csa_tree_add_14_36_groupi_n_2013 ();
drwire csa_tree_add_14_36_groupi_n_2014 ();
drwire csa_tree_add_14_36_groupi_n_2015 ();
drwire csa_tree_add_14_36_groupi_n_2016 ();
drwire csa_tree_add_14_36_groupi_n_2017 ();
drwire csa_tree_add_14_36_groupi_n_2018 ();
drwire csa_tree_add_14_36_groupi_n_2019 ();
drwire csa_tree_add_14_36_groupi_n_202 ();
drwire csa_tree_add_14_36_groupi_n_2020 ();
drwire csa_tree_add_14_36_groupi_n_2021 ();
drwire csa_tree_add_14_36_groupi_n_2022 ();
drwire csa_tree_add_14_36_groupi_n_2023 ();
drwire csa_tree_add_14_36_groupi_n_2024 ();
drwire csa_tree_add_14_36_groupi_n_2025 ();
drwire csa_tree_add_14_36_groupi_n_2026 ();
drwire csa_tree_add_14_36_groupi_n_2027 ();
drwire csa_tree_add_14_36_groupi_n_2028 ();
drwire csa_tree_add_14_36_groupi_n_2029 ();
drwire csa_tree_add_14_36_groupi_n_203 ();
drwire csa_tree_add_14_36_groupi_n_2030 ();
drwire csa_tree_add_14_36_groupi_n_2031 ();
drwire csa_tree_add_14_36_groupi_n_2032 ();
drwire csa_tree_add_14_36_groupi_n_2033 ();
drwire csa_tree_add_14_36_groupi_n_2034 ();
drwire csa_tree_add_14_36_groupi_n_2035 ();
drwire csa_tree_add_14_36_groupi_n_2036 ();
drwire csa_tree_add_14_36_groupi_n_2037 ();
drwire csa_tree_add_14_36_groupi_n_2038 ();
drwire csa_tree_add_14_36_groupi_n_2039 ();
drwire csa_tree_add_14_36_groupi_n_204 ();
drwire csa_tree_add_14_36_groupi_n_2040 ();
drwire csa_tree_add_14_36_groupi_n_2041 ();
drwire csa_tree_add_14_36_groupi_n_2042 ();
drwire csa_tree_add_14_36_groupi_n_2043 ();
drwire csa_tree_add_14_36_groupi_n_2044 ();
drwire csa_tree_add_14_36_groupi_n_2045 ();
drwire csa_tree_add_14_36_groupi_n_2046 ();
drwire csa_tree_add_14_36_groupi_n_2047 ();
drwire csa_tree_add_14_36_groupi_n_2048 ();
drwire csa_tree_add_14_36_groupi_n_2049 ();
drwire csa_tree_add_14_36_groupi_n_205 ();
drwire csa_tree_add_14_36_groupi_n_2050 ();
drwire csa_tree_add_14_36_groupi_n_2051 ();
drwire csa_tree_add_14_36_groupi_n_2052 ();
drwire csa_tree_add_14_36_groupi_n_2053 ();
drwire csa_tree_add_14_36_groupi_n_2054 ();
drwire csa_tree_add_14_36_groupi_n_2055 ();
drwire csa_tree_add_14_36_groupi_n_2056 ();
drwire csa_tree_add_14_36_groupi_n_2057 ();
drwire csa_tree_add_14_36_groupi_n_2058 ();
drwire csa_tree_add_14_36_groupi_n_2059 ();
drwire csa_tree_add_14_36_groupi_n_206 ();
drwire csa_tree_add_14_36_groupi_n_2060 ();
drwire csa_tree_add_14_36_groupi_n_2061 ();
drwire csa_tree_add_14_36_groupi_n_2062 ();
drwire csa_tree_add_14_36_groupi_n_2063 ();
drwire csa_tree_add_14_36_groupi_n_2064 ();
drwire csa_tree_add_14_36_groupi_n_2065 ();
drwire csa_tree_add_14_36_groupi_n_2066 ();
drwire csa_tree_add_14_36_groupi_n_2067 ();
drwire csa_tree_add_14_36_groupi_n_2068 ();
drwire csa_tree_add_14_36_groupi_n_2069 ();
drwire csa_tree_add_14_36_groupi_n_207 ();
drwire csa_tree_add_14_36_groupi_n_2070 ();
drwire csa_tree_add_14_36_groupi_n_2071 ();
drwire csa_tree_add_14_36_groupi_n_2072 ();
drwire csa_tree_add_14_36_groupi_n_2073 ();
drwire csa_tree_add_14_36_groupi_n_2074 ();
drwire csa_tree_add_14_36_groupi_n_2075 ();
drwire csa_tree_add_14_36_groupi_n_2076 ();
drwire csa_tree_add_14_36_groupi_n_2077 ();
drwire csa_tree_add_14_36_groupi_n_2078 ();
drwire csa_tree_add_14_36_groupi_n_2079 ();
drwire csa_tree_add_14_36_groupi_n_208 ();
drwire csa_tree_add_14_36_groupi_n_2080 ();
drwire csa_tree_add_14_36_groupi_n_2081 ();
drwire csa_tree_add_14_36_groupi_n_2082 ();
drwire csa_tree_add_14_36_groupi_n_2083 ();
drwire csa_tree_add_14_36_groupi_n_2084 ();
drwire csa_tree_add_14_36_groupi_n_2085 ();
drwire csa_tree_add_14_36_groupi_n_2086 ();
drwire csa_tree_add_14_36_groupi_n_2087 ();
drwire csa_tree_add_14_36_groupi_n_2088 ();
drwire csa_tree_add_14_36_groupi_n_2089 ();
drwire csa_tree_add_14_36_groupi_n_209 ();
drwire csa_tree_add_14_36_groupi_n_2090 ();
drwire csa_tree_add_14_36_groupi_n_2091 ();
drwire csa_tree_add_14_36_groupi_n_2092 ();
drwire csa_tree_add_14_36_groupi_n_2093 ();
drwire csa_tree_add_14_36_groupi_n_2094 ();
drwire csa_tree_add_14_36_groupi_n_2095 ();
drwire csa_tree_add_14_36_groupi_n_2096 ();
drwire csa_tree_add_14_36_groupi_n_2097 ();
drwire csa_tree_add_14_36_groupi_n_2098 ();
drwire csa_tree_add_14_36_groupi_n_2099 ();
drwire csa_tree_add_14_36_groupi_n_21 ();
drwire csa_tree_add_14_36_groupi_n_210 ();
drwire csa_tree_add_14_36_groupi_n_2100 ();
drwire csa_tree_add_14_36_groupi_n_2101 ();
drwire csa_tree_add_14_36_groupi_n_2102 ();
drwire csa_tree_add_14_36_groupi_n_2103 ();
drwire csa_tree_add_14_36_groupi_n_2104 ();
drwire csa_tree_add_14_36_groupi_n_2105 ();
drwire csa_tree_add_14_36_groupi_n_2106 ();
drwire csa_tree_add_14_36_groupi_n_2107 ();
drwire csa_tree_add_14_36_groupi_n_2108 ();
drwire csa_tree_add_14_36_groupi_n_2109 ();
drwire csa_tree_add_14_36_groupi_n_211 ();
drwire csa_tree_add_14_36_groupi_n_2110 ();
drwire csa_tree_add_14_36_groupi_n_2111 ();
drwire csa_tree_add_14_36_groupi_n_2112 ();
drwire csa_tree_add_14_36_groupi_n_2113 ();
drwire csa_tree_add_14_36_groupi_n_2114 ();
drwire csa_tree_add_14_36_groupi_n_2115 ();
drwire csa_tree_add_14_36_groupi_n_2116 ();
drwire csa_tree_add_14_36_groupi_n_2117 ();
drwire csa_tree_add_14_36_groupi_n_2118 ();
drwire csa_tree_add_14_36_groupi_n_2119 ();
drwire csa_tree_add_14_36_groupi_n_212 ();
drwire csa_tree_add_14_36_groupi_n_2120 ();
drwire csa_tree_add_14_36_groupi_n_2121 ();
drwire csa_tree_add_14_36_groupi_n_2122 ();
drwire csa_tree_add_14_36_groupi_n_2123 ();
drwire csa_tree_add_14_36_groupi_n_2124 ();
drwire csa_tree_add_14_36_groupi_n_2125 ();
drwire csa_tree_add_14_36_groupi_n_2126 ();
drwire csa_tree_add_14_36_groupi_n_2127 ();
drwire csa_tree_add_14_36_groupi_n_2128 ();
drwire csa_tree_add_14_36_groupi_n_2129 ();
drwire csa_tree_add_14_36_groupi_n_213 ();
drwire csa_tree_add_14_36_groupi_n_2130 ();
drwire csa_tree_add_14_36_groupi_n_2131 ();
drwire csa_tree_add_14_36_groupi_n_2132 ();
drwire csa_tree_add_14_36_groupi_n_2133 ();
drwire csa_tree_add_14_36_groupi_n_2134 ();
drwire csa_tree_add_14_36_groupi_n_2135 ();
drwire csa_tree_add_14_36_groupi_n_2136 ();
drwire csa_tree_add_14_36_groupi_n_2137 ();
drwire csa_tree_add_14_36_groupi_n_2138 ();
drwire csa_tree_add_14_36_groupi_n_2139 ();
drwire csa_tree_add_14_36_groupi_n_214 ();
drwire csa_tree_add_14_36_groupi_n_2140 ();
drwire csa_tree_add_14_36_groupi_n_2141 ();
drwire csa_tree_add_14_36_groupi_n_2142 ();
drwire csa_tree_add_14_36_groupi_n_2143 ();
drwire csa_tree_add_14_36_groupi_n_2144 ();
drwire csa_tree_add_14_36_groupi_n_2145 ();
drwire csa_tree_add_14_36_groupi_n_2146 ();
drwire csa_tree_add_14_36_groupi_n_2147 ();
drwire csa_tree_add_14_36_groupi_n_2148 ();
drwire csa_tree_add_14_36_groupi_n_2149 ();
drwire csa_tree_add_14_36_groupi_n_215 ();
drwire csa_tree_add_14_36_groupi_n_2150 ();
drwire csa_tree_add_14_36_groupi_n_2151 ();
drwire csa_tree_add_14_36_groupi_n_2152 ();
drwire csa_tree_add_14_36_groupi_n_2153 ();
drwire csa_tree_add_14_36_groupi_n_2154 ();
drwire csa_tree_add_14_36_groupi_n_2155 ();
drwire csa_tree_add_14_36_groupi_n_2156 ();
drwire csa_tree_add_14_36_groupi_n_2157 ();
drwire csa_tree_add_14_36_groupi_n_2158 ();
drwire csa_tree_add_14_36_groupi_n_2159 ();
drwire csa_tree_add_14_36_groupi_n_216 ();
drwire csa_tree_add_14_36_groupi_n_2160 ();
drwire csa_tree_add_14_36_groupi_n_2161 ();
drwire csa_tree_add_14_36_groupi_n_2162 ();
drwire csa_tree_add_14_36_groupi_n_2163 ();
drwire csa_tree_add_14_36_groupi_n_2164 ();
drwire csa_tree_add_14_36_groupi_n_2165 ();
drwire csa_tree_add_14_36_groupi_n_2166 ();
drwire csa_tree_add_14_36_groupi_n_2167 ();
drwire csa_tree_add_14_36_groupi_n_2168 ();
drwire csa_tree_add_14_36_groupi_n_2169 ();
drwire csa_tree_add_14_36_groupi_n_217 ();
drwire csa_tree_add_14_36_groupi_n_2170 ();
drwire csa_tree_add_14_36_groupi_n_2171 ();
drwire csa_tree_add_14_36_groupi_n_2172 ();
drwire csa_tree_add_14_36_groupi_n_2173 ();
drwire csa_tree_add_14_36_groupi_n_2174 ();
drwire csa_tree_add_14_36_groupi_n_2175 ();
drwire csa_tree_add_14_36_groupi_n_2176 ();
drwire csa_tree_add_14_36_groupi_n_2177 ();
drwire csa_tree_add_14_36_groupi_n_2178 ();
drwire csa_tree_add_14_36_groupi_n_2179 ();
drwire csa_tree_add_14_36_groupi_n_218 ();
drwire csa_tree_add_14_36_groupi_n_2180 ();
drwire csa_tree_add_14_36_groupi_n_2181 ();
drwire csa_tree_add_14_36_groupi_n_2182 ();
drwire csa_tree_add_14_36_groupi_n_2183 ();
drwire csa_tree_add_14_36_groupi_n_2184 ();
drwire csa_tree_add_14_36_groupi_n_2185 ();
drwire csa_tree_add_14_36_groupi_n_2186 ();
drwire csa_tree_add_14_36_groupi_n_2187 ();
drwire csa_tree_add_14_36_groupi_n_2188 ();
drwire csa_tree_add_14_36_groupi_n_2189 ();
drwire csa_tree_add_14_36_groupi_n_219 ();
drwire csa_tree_add_14_36_groupi_n_2190 ();
drwire csa_tree_add_14_36_groupi_n_2191 ();
drwire csa_tree_add_14_36_groupi_n_2192 ();
drwire csa_tree_add_14_36_groupi_n_2193 ();
drwire csa_tree_add_14_36_groupi_n_2194 ();
drwire csa_tree_add_14_36_groupi_n_2195 ();
drwire csa_tree_add_14_36_groupi_n_2196 ();
drwire csa_tree_add_14_36_groupi_n_2197 ();
drwire csa_tree_add_14_36_groupi_n_2198 ();
drwire csa_tree_add_14_36_groupi_n_2199 ();
drwire csa_tree_add_14_36_groupi_n_220 ();
drwire csa_tree_add_14_36_groupi_n_2200 ();
drwire csa_tree_add_14_36_groupi_n_2201 ();
drwire csa_tree_add_14_36_groupi_n_2202 ();
drwire csa_tree_add_14_36_groupi_n_2203 ();
drwire csa_tree_add_14_36_groupi_n_2204 ();
drwire csa_tree_add_14_36_groupi_n_2205 ();
drwire csa_tree_add_14_36_groupi_n_2206 ();
drwire csa_tree_add_14_36_groupi_n_2207 ();
drwire csa_tree_add_14_36_groupi_n_2208 ();
drwire csa_tree_add_14_36_groupi_n_2209 ();
drwire csa_tree_add_14_36_groupi_n_221 ();
drwire csa_tree_add_14_36_groupi_n_2210 ();
drwire csa_tree_add_14_36_groupi_n_2211 ();
drwire csa_tree_add_14_36_groupi_n_2212 ();
drwire csa_tree_add_14_36_groupi_n_2213 ();
drwire csa_tree_add_14_36_groupi_n_2214 ();
drwire csa_tree_add_14_36_groupi_n_2215 ();
drwire csa_tree_add_14_36_groupi_n_2216 ();
drwire csa_tree_add_14_36_groupi_n_2217 ();
drwire csa_tree_add_14_36_groupi_n_2218 ();
drwire csa_tree_add_14_36_groupi_n_2219 ();
drwire csa_tree_add_14_36_groupi_n_222 ();
drwire csa_tree_add_14_36_groupi_n_2220 ();
drwire csa_tree_add_14_36_groupi_n_2221 ();
drwire csa_tree_add_14_36_groupi_n_2222 ();
drwire csa_tree_add_14_36_groupi_n_2223 ();
drwire csa_tree_add_14_36_groupi_n_2224 ();
drwire csa_tree_add_14_36_groupi_n_2225 ();
drwire csa_tree_add_14_36_groupi_n_2226 ();
drwire csa_tree_add_14_36_groupi_n_2227 ();
drwire csa_tree_add_14_36_groupi_n_2228 ();
drwire csa_tree_add_14_36_groupi_n_2229 ();
drwire csa_tree_add_14_36_groupi_n_223 ();
drwire csa_tree_add_14_36_groupi_n_2230 ();
drwire csa_tree_add_14_36_groupi_n_2231 ();
drwire csa_tree_add_14_36_groupi_n_2232 ();
drwire csa_tree_add_14_36_groupi_n_2233 ();
drwire csa_tree_add_14_36_groupi_n_2234 ();
drwire csa_tree_add_14_36_groupi_n_2235 ();
drwire csa_tree_add_14_36_groupi_n_2236 ();
drwire csa_tree_add_14_36_groupi_n_2237 ();
drwire csa_tree_add_14_36_groupi_n_2238 ();
drwire csa_tree_add_14_36_groupi_n_2239 ();
drwire csa_tree_add_14_36_groupi_n_224 ();
drwire csa_tree_add_14_36_groupi_n_2240 ();
drwire csa_tree_add_14_36_groupi_n_2241 ();
drwire csa_tree_add_14_36_groupi_n_2242 ();
drwire csa_tree_add_14_36_groupi_n_2243 ();
drwire csa_tree_add_14_36_groupi_n_2244 ();
drwire csa_tree_add_14_36_groupi_n_2245 ();
drwire csa_tree_add_14_36_groupi_n_2246 ();
drwire csa_tree_add_14_36_groupi_n_2247 ();
drwire csa_tree_add_14_36_groupi_n_2248 ();
drwire csa_tree_add_14_36_groupi_n_2249 ();
drwire csa_tree_add_14_36_groupi_n_225 ();
drwire csa_tree_add_14_36_groupi_n_2250 ();
drwire csa_tree_add_14_36_groupi_n_2251 ();
drwire csa_tree_add_14_36_groupi_n_2252 ();
drwire csa_tree_add_14_36_groupi_n_2253 ();
drwire csa_tree_add_14_36_groupi_n_2254 ();
drwire csa_tree_add_14_36_groupi_n_2255 ();
drwire csa_tree_add_14_36_groupi_n_2256 ();
drwire csa_tree_add_14_36_groupi_n_2257 ();
drwire csa_tree_add_14_36_groupi_n_2258 ();
drwire csa_tree_add_14_36_groupi_n_2259 ();
drwire csa_tree_add_14_36_groupi_n_226 ();
drwire csa_tree_add_14_36_groupi_n_2260 ();
drwire csa_tree_add_14_36_groupi_n_2261 ();
drwire csa_tree_add_14_36_groupi_n_2262 ();
drwire csa_tree_add_14_36_groupi_n_2263 ();
drwire csa_tree_add_14_36_groupi_n_2264 ();
drwire csa_tree_add_14_36_groupi_n_2265 ();
drwire csa_tree_add_14_36_groupi_n_2266 ();
drwire csa_tree_add_14_36_groupi_n_2267 ();
drwire csa_tree_add_14_36_groupi_n_2268 ();
drwire csa_tree_add_14_36_groupi_n_2269 ();
drwire csa_tree_add_14_36_groupi_n_227 ();
drwire csa_tree_add_14_36_groupi_n_2270 ();
drwire csa_tree_add_14_36_groupi_n_2271 ();
drwire csa_tree_add_14_36_groupi_n_2272 ();
drwire csa_tree_add_14_36_groupi_n_2275 ();
drwire csa_tree_add_14_36_groupi_n_2276 ();
drwire csa_tree_add_14_36_groupi_n_2277 ();
drwire csa_tree_add_14_36_groupi_n_2278 ();
drwire csa_tree_add_14_36_groupi_n_2279 ();
drwire csa_tree_add_14_36_groupi_n_228 ();
drwire csa_tree_add_14_36_groupi_n_2280 ();
drwire csa_tree_add_14_36_groupi_n_2281 ();
drwire csa_tree_add_14_36_groupi_n_2282 ();
drwire csa_tree_add_14_36_groupi_n_2283 ();
drwire csa_tree_add_14_36_groupi_n_2284 ();
drwire csa_tree_add_14_36_groupi_n_2285 ();
drwire csa_tree_add_14_36_groupi_n_2286 ();
drwire csa_tree_add_14_36_groupi_n_2287 ();
drwire csa_tree_add_14_36_groupi_n_2288 ();
drwire csa_tree_add_14_36_groupi_n_2291 ();
drwire csa_tree_add_14_36_groupi_n_2292 ();
drwire csa_tree_add_14_36_groupi_n_2293 ();
drwire csa_tree_add_14_36_groupi_n_2294 ();
drwire csa_tree_add_14_36_groupi_n_2295 ();
drwire csa_tree_add_14_36_groupi_n_2297 ();
drwire csa_tree_add_14_36_groupi_n_2298 ();
drwire csa_tree_add_14_36_groupi_n_2299 ();
drwire csa_tree_add_14_36_groupi_n_23 ();
drwire csa_tree_add_14_36_groupi_n_230 ();
drwire csa_tree_add_14_36_groupi_n_2300 ();
drwire csa_tree_add_14_36_groupi_n_2301 ();
drwire csa_tree_add_14_36_groupi_n_2302 ();
drwire csa_tree_add_14_36_groupi_n_2303 ();
drwire csa_tree_add_14_36_groupi_n_2304 ();
drwire csa_tree_add_14_36_groupi_n_2305 ();
drwire csa_tree_add_14_36_groupi_n_2306 ();
drwire csa_tree_add_14_36_groupi_n_2307 ();
drwire csa_tree_add_14_36_groupi_n_2308 ();
drwire csa_tree_add_14_36_groupi_n_2309 ();
drwire csa_tree_add_14_36_groupi_n_231 ();
drwire csa_tree_add_14_36_groupi_n_2310 ();
drwire csa_tree_add_14_36_groupi_n_2311 ();
drwire csa_tree_add_14_36_groupi_n_2312 ();
drwire csa_tree_add_14_36_groupi_n_2313 ();
drwire csa_tree_add_14_36_groupi_n_2314 ();
drwire csa_tree_add_14_36_groupi_n_2315 ();
drwire csa_tree_add_14_36_groupi_n_2316 ();
drwire csa_tree_add_14_36_groupi_n_2317 ();
drwire csa_tree_add_14_36_groupi_n_2318 ();
drwire csa_tree_add_14_36_groupi_n_2319 ();
drwire csa_tree_add_14_36_groupi_n_2320 ();
drwire csa_tree_add_14_36_groupi_n_2321 ();
drwire csa_tree_add_14_36_groupi_n_234 ();
drwire csa_tree_add_14_36_groupi_n_235 ();
drwire csa_tree_add_14_36_groupi_n_236 ();
drwire csa_tree_add_14_36_groupi_n_237 ();
drwire csa_tree_add_14_36_groupi_n_238 ();
drwire csa_tree_add_14_36_groupi_n_239 ();
drwire csa_tree_add_14_36_groupi_n_24 ();
drwire csa_tree_add_14_36_groupi_n_240 ();
drwire csa_tree_add_14_36_groupi_n_241 ();
drwire csa_tree_add_14_36_groupi_n_2410 ();
drwire csa_tree_add_14_36_groupi_n_2412 ();
drwire csa_tree_add_14_36_groupi_n_2416 ();
drwire csa_tree_add_14_36_groupi_n_242 ();
drwire csa_tree_add_14_36_groupi_n_243 ();
drwire csa_tree_add_14_36_groupi_n_245 ();
drwire csa_tree_add_14_36_groupi_n_246 ();
drwire csa_tree_add_14_36_groupi_n_247 ();
drwire csa_tree_add_14_36_groupi_n_248 ();
drwire csa_tree_add_14_36_groupi_n_249 ();
drwire csa_tree_add_14_36_groupi_n_25 ();
drwire csa_tree_add_14_36_groupi_n_250 ();
drwire csa_tree_add_14_36_groupi_n_251 ();
drwire csa_tree_add_14_36_groupi_n_252 ();
drwire csa_tree_add_14_36_groupi_n_253 ();
drwire csa_tree_add_14_36_groupi_n_254 ();
drwire csa_tree_add_14_36_groupi_n_255 ();
drwire csa_tree_add_14_36_groupi_n_257 ();
drwire csa_tree_add_14_36_groupi_n_259 ();
drwire csa_tree_add_14_36_groupi_n_26 ();
drwire csa_tree_add_14_36_groupi_n_260 ();
drwire csa_tree_add_14_36_groupi_n_261 ();
drwire csa_tree_add_14_36_groupi_n_262 ();
drwire csa_tree_add_14_36_groupi_n_263 ();
drwire csa_tree_add_14_36_groupi_n_264 ();
drwire csa_tree_add_14_36_groupi_n_265 ();
drwire csa_tree_add_14_36_groupi_n_266 ();
drwire csa_tree_add_14_36_groupi_n_267 ();
drwire csa_tree_add_14_36_groupi_n_268 ();
drwire csa_tree_add_14_36_groupi_n_269 ();
drwire csa_tree_add_14_36_groupi_n_27 ();
drwire csa_tree_add_14_36_groupi_n_270 ();
drwire csa_tree_add_14_36_groupi_n_271 ();
drwire csa_tree_add_14_36_groupi_n_272 ();
drwire csa_tree_add_14_36_groupi_n_273 ();
drwire csa_tree_add_14_36_groupi_n_274 ();
drwire csa_tree_add_14_36_groupi_n_275 ();
drwire csa_tree_add_14_36_groupi_n_276 ();
drwire csa_tree_add_14_36_groupi_n_277 ();
drwire csa_tree_add_14_36_groupi_n_278 ();
drwire csa_tree_add_14_36_groupi_n_279 ();
drwire csa_tree_add_14_36_groupi_n_28 ();
drwire csa_tree_add_14_36_groupi_n_280 ();
drwire csa_tree_add_14_36_groupi_n_281 ();
drwire csa_tree_add_14_36_groupi_n_282 ();
drwire csa_tree_add_14_36_groupi_n_283 ();
drwire csa_tree_add_14_36_groupi_n_284 ();
drwire csa_tree_add_14_36_groupi_n_285 ();
drwire csa_tree_add_14_36_groupi_n_286 ();
drwire csa_tree_add_14_36_groupi_n_287 ();
drwire csa_tree_add_14_36_groupi_n_288 ();
drwire csa_tree_add_14_36_groupi_n_289 ();
drwire csa_tree_add_14_36_groupi_n_29 ();
drwire csa_tree_add_14_36_groupi_n_290 ();
drwire csa_tree_add_14_36_groupi_n_291 ();
drwire csa_tree_add_14_36_groupi_n_292 ();
drwire csa_tree_add_14_36_groupi_n_293 ();
drwire csa_tree_add_14_36_groupi_n_294 ();
drwire csa_tree_add_14_36_groupi_n_295 ();
drwire csa_tree_add_14_36_groupi_n_296 ();
drwire csa_tree_add_14_36_groupi_n_297 ();
drwire csa_tree_add_14_36_groupi_n_298 ();
drwire csa_tree_add_14_36_groupi_n_299 ();
drwire csa_tree_add_14_36_groupi_n_3 ();
drwire csa_tree_add_14_36_groupi_n_30 ();
drwire csa_tree_add_14_36_groupi_n_300 ();
drwire csa_tree_add_14_36_groupi_n_301 ();
drwire csa_tree_add_14_36_groupi_n_302 ();
drwire csa_tree_add_14_36_groupi_n_303 ();
drwire csa_tree_add_14_36_groupi_n_304 ();
drwire csa_tree_add_14_36_groupi_n_305 ();
drwire csa_tree_add_14_36_groupi_n_306 ();
drwire csa_tree_add_14_36_groupi_n_307 ();
drwire csa_tree_add_14_36_groupi_n_308 ();
drwire csa_tree_add_14_36_groupi_n_309 ();
drwire csa_tree_add_14_36_groupi_n_31 ();
drwire csa_tree_add_14_36_groupi_n_310 ();
drwire csa_tree_add_14_36_groupi_n_311 ();
drwire csa_tree_add_14_36_groupi_n_312 ();
drwire csa_tree_add_14_36_groupi_n_313 ();
drwire csa_tree_add_14_36_groupi_n_315 ();
drwire csa_tree_add_14_36_groupi_n_316 ();
drwire csa_tree_add_14_36_groupi_n_317 ();
drwire csa_tree_add_14_36_groupi_n_318 ();
drwire csa_tree_add_14_36_groupi_n_319 ();
drwire csa_tree_add_14_36_groupi_n_32 ();
drwire csa_tree_add_14_36_groupi_n_320 ();
drwire csa_tree_add_14_36_groupi_n_321 ();
drwire csa_tree_add_14_36_groupi_n_322 ();
drwire csa_tree_add_14_36_groupi_n_323 ();
drwire csa_tree_add_14_36_groupi_n_324 ();
drwire csa_tree_add_14_36_groupi_n_325 ();
drwire csa_tree_add_14_36_groupi_n_326 ();
drwire csa_tree_add_14_36_groupi_n_327 ();
drwire csa_tree_add_14_36_groupi_n_328 ();
drwire csa_tree_add_14_36_groupi_n_329 ();
drwire csa_tree_add_14_36_groupi_n_33 ();
drwire csa_tree_add_14_36_groupi_n_330 ();
drwire csa_tree_add_14_36_groupi_n_331 ();
drwire csa_tree_add_14_36_groupi_n_332 ();
drwire csa_tree_add_14_36_groupi_n_333 ();
drwire csa_tree_add_14_36_groupi_n_334 ();
drwire csa_tree_add_14_36_groupi_n_335 ();
drwire csa_tree_add_14_36_groupi_n_336 ();
drwire csa_tree_add_14_36_groupi_n_337 ();
drwire csa_tree_add_14_36_groupi_n_338 ();
drwire csa_tree_add_14_36_groupi_n_339 ();
drwire csa_tree_add_14_36_groupi_n_34 ();
drwire csa_tree_add_14_36_groupi_n_340 ();
drwire csa_tree_add_14_36_groupi_n_341 ();
drwire csa_tree_add_14_36_groupi_n_342 ();
drwire csa_tree_add_14_36_groupi_n_343 ();
drwire csa_tree_add_14_36_groupi_n_344 ();
drwire csa_tree_add_14_36_groupi_n_345 ();
drwire csa_tree_add_14_36_groupi_n_346 ();
drwire csa_tree_add_14_36_groupi_n_347 ();
drwire csa_tree_add_14_36_groupi_n_348 ();
drwire csa_tree_add_14_36_groupi_n_349 ();
drwire csa_tree_add_14_36_groupi_n_35 ();
drwire csa_tree_add_14_36_groupi_n_350 ();
drwire csa_tree_add_14_36_groupi_n_351 ();
drwire csa_tree_add_14_36_groupi_n_352 ();
drwire csa_tree_add_14_36_groupi_n_353 ();
drwire csa_tree_add_14_36_groupi_n_354 ();
drwire csa_tree_add_14_36_groupi_n_355 ();
drwire csa_tree_add_14_36_groupi_n_356 ();
drwire csa_tree_add_14_36_groupi_n_357 ();
drwire csa_tree_add_14_36_groupi_n_358 ();
drwire csa_tree_add_14_36_groupi_n_359 ();
drwire csa_tree_add_14_36_groupi_n_36 ();
drwire csa_tree_add_14_36_groupi_n_360 ();
drwire csa_tree_add_14_36_groupi_n_361 ();
drwire csa_tree_add_14_36_groupi_n_362 ();
drwire csa_tree_add_14_36_groupi_n_363 ();
drwire csa_tree_add_14_36_groupi_n_364 ();
drwire csa_tree_add_14_36_groupi_n_365 ();
drwire csa_tree_add_14_36_groupi_n_366 ();
drwire csa_tree_add_14_36_groupi_n_367 ();
drwire csa_tree_add_14_36_groupi_n_368 ();
drwire csa_tree_add_14_36_groupi_n_369 ();
drwire csa_tree_add_14_36_groupi_n_37 ();
drwire csa_tree_add_14_36_groupi_n_370 ();
drwire csa_tree_add_14_36_groupi_n_371 ();
drwire csa_tree_add_14_36_groupi_n_372 ();
drwire csa_tree_add_14_36_groupi_n_373 ();
drwire csa_tree_add_14_36_groupi_n_374 ();
drwire csa_tree_add_14_36_groupi_n_375 ();
drwire csa_tree_add_14_36_groupi_n_376 ();
drwire csa_tree_add_14_36_groupi_n_377 ();
drwire csa_tree_add_14_36_groupi_n_378 ();
drwire csa_tree_add_14_36_groupi_n_379 ();
drwire csa_tree_add_14_36_groupi_n_38 ();
drwire csa_tree_add_14_36_groupi_n_380 ();
drwire csa_tree_add_14_36_groupi_n_381 ();
drwire csa_tree_add_14_36_groupi_n_382 ();
drwire csa_tree_add_14_36_groupi_n_383 ();
drwire csa_tree_add_14_36_groupi_n_384 ();
drwire csa_tree_add_14_36_groupi_n_385 ();
drwire csa_tree_add_14_36_groupi_n_386 ();
drwire csa_tree_add_14_36_groupi_n_387 ();
drwire csa_tree_add_14_36_groupi_n_388 ();
drwire csa_tree_add_14_36_groupi_n_389 ();
drwire csa_tree_add_14_36_groupi_n_39 ();
drwire csa_tree_add_14_36_groupi_n_390 ();
drwire csa_tree_add_14_36_groupi_n_391 ();
drwire csa_tree_add_14_36_groupi_n_392 ();
drwire csa_tree_add_14_36_groupi_n_393 ();
drwire csa_tree_add_14_36_groupi_n_395 ();
drwire csa_tree_add_14_36_groupi_n_397 ();
drwire csa_tree_add_14_36_groupi_n_399 ();
drwire csa_tree_add_14_36_groupi_n_4 ();
drwire csa_tree_add_14_36_groupi_n_40 ();
drwire csa_tree_add_14_36_groupi_n_401 ();
drwire csa_tree_add_14_36_groupi_n_403 ();
drwire csa_tree_add_14_36_groupi_n_404 ();
drwire csa_tree_add_14_36_groupi_n_405 ();
drwire csa_tree_add_14_36_groupi_n_406 ();
drwire csa_tree_add_14_36_groupi_n_407 ();
drwire csa_tree_add_14_36_groupi_n_408 ();
drwire csa_tree_add_14_36_groupi_n_409 ();
drwire csa_tree_add_14_36_groupi_n_41 ();
drwire csa_tree_add_14_36_groupi_n_410 ();
drwire csa_tree_add_14_36_groupi_n_411 ();
drwire csa_tree_add_14_36_groupi_n_412 ();
drwire csa_tree_add_14_36_groupi_n_413 ();
drwire csa_tree_add_14_36_groupi_n_414 ();
drwire csa_tree_add_14_36_groupi_n_415 ();
drwire csa_tree_add_14_36_groupi_n_416 ();
drwire csa_tree_add_14_36_groupi_n_417 ();
drwire csa_tree_add_14_36_groupi_n_418 ();
drwire csa_tree_add_14_36_groupi_n_419 ();
drwire csa_tree_add_14_36_groupi_n_42 ();
drwire csa_tree_add_14_36_groupi_n_420 ();
drwire csa_tree_add_14_36_groupi_n_421 ();
drwire csa_tree_add_14_36_groupi_n_422 ();
drwire csa_tree_add_14_36_groupi_n_423 ();
drwire csa_tree_add_14_36_groupi_n_424 ();
drwire csa_tree_add_14_36_groupi_n_425 ();
drwire csa_tree_add_14_36_groupi_n_426 ();
drwire csa_tree_add_14_36_groupi_n_427 ();
drwire csa_tree_add_14_36_groupi_n_428 ();
drwire csa_tree_add_14_36_groupi_n_429 ();
drwire csa_tree_add_14_36_groupi_n_43 ();
drwire csa_tree_add_14_36_groupi_n_430 ();
drwire csa_tree_add_14_36_groupi_n_431 ();
drwire csa_tree_add_14_36_groupi_n_432 ();
drwire csa_tree_add_14_36_groupi_n_433 ();
drwire csa_tree_add_14_36_groupi_n_434 ();
drwire csa_tree_add_14_36_groupi_n_435 ();
drwire csa_tree_add_14_36_groupi_n_436 ();
drwire csa_tree_add_14_36_groupi_n_437 ();
drwire csa_tree_add_14_36_groupi_n_438 ();
drwire csa_tree_add_14_36_groupi_n_439 ();
drwire csa_tree_add_14_36_groupi_n_44 ();
drwire csa_tree_add_14_36_groupi_n_440 ();
drwire csa_tree_add_14_36_groupi_n_441 ();
drwire csa_tree_add_14_36_groupi_n_442 ();
drwire csa_tree_add_14_36_groupi_n_443 ();
drwire csa_tree_add_14_36_groupi_n_444 ();
drwire csa_tree_add_14_36_groupi_n_445 ();
drwire csa_tree_add_14_36_groupi_n_446 ();
drwire csa_tree_add_14_36_groupi_n_447 ();
drwire csa_tree_add_14_36_groupi_n_448 ();
drwire csa_tree_add_14_36_groupi_n_449 ();
drwire csa_tree_add_14_36_groupi_n_45 ();
drwire csa_tree_add_14_36_groupi_n_450 ();
drwire csa_tree_add_14_36_groupi_n_451 ();
drwire csa_tree_add_14_36_groupi_n_452 ();
drwire csa_tree_add_14_36_groupi_n_453 ();
drwire csa_tree_add_14_36_groupi_n_454 ();
drwire csa_tree_add_14_36_groupi_n_455 ();
drwire csa_tree_add_14_36_groupi_n_456 ();
drwire csa_tree_add_14_36_groupi_n_457 ();
drwire csa_tree_add_14_36_groupi_n_458 ();
drwire csa_tree_add_14_36_groupi_n_459 ();
drwire csa_tree_add_14_36_groupi_n_46 ();
drwire csa_tree_add_14_36_groupi_n_460 ();
drwire csa_tree_add_14_36_groupi_n_461 ();
drwire csa_tree_add_14_36_groupi_n_462 ();
drwire csa_tree_add_14_36_groupi_n_463 ();
drwire csa_tree_add_14_36_groupi_n_464 ();
drwire csa_tree_add_14_36_groupi_n_465 ();
drwire csa_tree_add_14_36_groupi_n_466 ();
drwire csa_tree_add_14_36_groupi_n_467 ();
drwire csa_tree_add_14_36_groupi_n_468 ();
drwire csa_tree_add_14_36_groupi_n_469 ();
drwire csa_tree_add_14_36_groupi_n_470 ();
drwire csa_tree_add_14_36_groupi_n_471 ();
drwire csa_tree_add_14_36_groupi_n_472 ();
drwire csa_tree_add_14_36_groupi_n_473 ();
drwire csa_tree_add_14_36_groupi_n_474 ();
drwire csa_tree_add_14_36_groupi_n_475 ();
drwire csa_tree_add_14_36_groupi_n_476 ();
drwire csa_tree_add_14_36_groupi_n_477 ();
drwire csa_tree_add_14_36_groupi_n_478 ();
drwire csa_tree_add_14_36_groupi_n_479 ();
drwire csa_tree_add_14_36_groupi_n_48 ();
drwire csa_tree_add_14_36_groupi_n_480 ();
drwire csa_tree_add_14_36_groupi_n_481 ();
drwire csa_tree_add_14_36_groupi_n_482 ();
drwire csa_tree_add_14_36_groupi_n_483 ();
drwire csa_tree_add_14_36_groupi_n_484 ();
drwire csa_tree_add_14_36_groupi_n_485 ();
drwire csa_tree_add_14_36_groupi_n_486 ();
drwire csa_tree_add_14_36_groupi_n_487 ();
drwire csa_tree_add_14_36_groupi_n_488 ();
drwire csa_tree_add_14_36_groupi_n_489 ();
drwire csa_tree_add_14_36_groupi_n_49 ();
drwire csa_tree_add_14_36_groupi_n_490 ();
drwire csa_tree_add_14_36_groupi_n_491 ();
drwire csa_tree_add_14_36_groupi_n_492 ();
drwire csa_tree_add_14_36_groupi_n_493 ();
drwire csa_tree_add_14_36_groupi_n_495 ();
drwire csa_tree_add_14_36_groupi_n_496 ();
drwire csa_tree_add_14_36_groupi_n_497 ();
drwire csa_tree_add_14_36_groupi_n_498 ();
drwire csa_tree_add_14_36_groupi_n_499 ();
drwire csa_tree_add_14_36_groupi_n_5 ();
drwire csa_tree_add_14_36_groupi_n_50 ();
drwire csa_tree_add_14_36_groupi_n_500 ();
drwire csa_tree_add_14_36_groupi_n_501 ();
drwire csa_tree_add_14_36_groupi_n_502 ();
drwire csa_tree_add_14_36_groupi_n_503 ();
drwire csa_tree_add_14_36_groupi_n_504 ();
drwire csa_tree_add_14_36_groupi_n_505 ();
drwire csa_tree_add_14_36_groupi_n_506 ();
drwire csa_tree_add_14_36_groupi_n_507 ();
drwire csa_tree_add_14_36_groupi_n_51 ();
drwire csa_tree_add_14_36_groupi_n_513 ();
drwire csa_tree_add_14_36_groupi_n_515 ();
drwire csa_tree_add_14_36_groupi_n_516 ();
drwire csa_tree_add_14_36_groupi_n_517 ();
drwire csa_tree_add_14_36_groupi_n_518 ();
drwire csa_tree_add_14_36_groupi_n_519 ();
drwire csa_tree_add_14_36_groupi_n_52 ();
drwire csa_tree_add_14_36_groupi_n_520 ();
drwire csa_tree_add_14_36_groupi_n_521 ();
drwire csa_tree_add_14_36_groupi_n_522 ();
drwire csa_tree_add_14_36_groupi_n_523 ();
drwire csa_tree_add_14_36_groupi_n_524 ();
drwire csa_tree_add_14_36_groupi_n_525 ();
drwire csa_tree_add_14_36_groupi_n_526 ();
drwire csa_tree_add_14_36_groupi_n_527 ();
drwire csa_tree_add_14_36_groupi_n_528 ();
drwire csa_tree_add_14_36_groupi_n_529 ();
drwire csa_tree_add_14_36_groupi_n_53 ();
drwire csa_tree_add_14_36_groupi_n_530 ();
drwire csa_tree_add_14_36_groupi_n_531 ();
drwire csa_tree_add_14_36_groupi_n_532 ();
drwire csa_tree_add_14_36_groupi_n_533 ();
drwire csa_tree_add_14_36_groupi_n_534 ();
drwire csa_tree_add_14_36_groupi_n_535 ();
drwire csa_tree_add_14_36_groupi_n_536 ();
drwire csa_tree_add_14_36_groupi_n_537 ();
drwire csa_tree_add_14_36_groupi_n_538 ();
drwire csa_tree_add_14_36_groupi_n_539 ();
drwire csa_tree_add_14_36_groupi_n_54 ();
drwire csa_tree_add_14_36_groupi_n_540 ();
drwire csa_tree_add_14_36_groupi_n_541 ();
drwire csa_tree_add_14_36_groupi_n_542 ();
drwire csa_tree_add_14_36_groupi_n_543 ();
drwire csa_tree_add_14_36_groupi_n_544 ();
drwire csa_tree_add_14_36_groupi_n_545 ();
drwire csa_tree_add_14_36_groupi_n_546 ();
drwire csa_tree_add_14_36_groupi_n_547 ();
drwire csa_tree_add_14_36_groupi_n_548 ();
drwire csa_tree_add_14_36_groupi_n_549 ();
drwire csa_tree_add_14_36_groupi_n_550 ();
drwire csa_tree_add_14_36_groupi_n_551 ();
drwire csa_tree_add_14_36_groupi_n_552 ();
drwire csa_tree_add_14_36_groupi_n_553 ();
drwire csa_tree_add_14_36_groupi_n_554 ();
drwire csa_tree_add_14_36_groupi_n_555 ();
drwire csa_tree_add_14_36_groupi_n_556 ();
drwire csa_tree_add_14_36_groupi_n_557 ();
drwire csa_tree_add_14_36_groupi_n_558 ();
drwire csa_tree_add_14_36_groupi_n_559 ();
drwire csa_tree_add_14_36_groupi_n_56 ();
drwire csa_tree_add_14_36_groupi_n_560 ();
drwire csa_tree_add_14_36_groupi_n_561 ();
drwire csa_tree_add_14_36_groupi_n_562 ();
drwire csa_tree_add_14_36_groupi_n_563 ();
drwire csa_tree_add_14_36_groupi_n_564 ();
drwire csa_tree_add_14_36_groupi_n_565 ();
drwire csa_tree_add_14_36_groupi_n_566 ();
drwire csa_tree_add_14_36_groupi_n_567 ();
drwire csa_tree_add_14_36_groupi_n_568 ();
drwire csa_tree_add_14_36_groupi_n_569 ();
drwire csa_tree_add_14_36_groupi_n_57 ();
drwire csa_tree_add_14_36_groupi_n_570 ();
drwire csa_tree_add_14_36_groupi_n_571 ();
drwire csa_tree_add_14_36_groupi_n_572 ();
drwire csa_tree_add_14_36_groupi_n_573 ();
drwire csa_tree_add_14_36_groupi_n_574 ();
drwire csa_tree_add_14_36_groupi_n_575 ();
drwire csa_tree_add_14_36_groupi_n_576 ();
drwire csa_tree_add_14_36_groupi_n_577 ();
drwire csa_tree_add_14_36_groupi_n_578 ();
drwire csa_tree_add_14_36_groupi_n_579 ();
drwire csa_tree_add_14_36_groupi_n_580 ();
drwire csa_tree_add_14_36_groupi_n_581 ();
drwire csa_tree_add_14_36_groupi_n_582 ();
drwire csa_tree_add_14_36_groupi_n_583 ();
drwire csa_tree_add_14_36_groupi_n_584 ();
drwire csa_tree_add_14_36_groupi_n_585 ();
drwire csa_tree_add_14_36_groupi_n_586 ();
drwire csa_tree_add_14_36_groupi_n_587 ();
drwire csa_tree_add_14_36_groupi_n_588 ();
drwire csa_tree_add_14_36_groupi_n_589 ();
drwire csa_tree_add_14_36_groupi_n_59 ();
drwire csa_tree_add_14_36_groupi_n_590 ();
drwire csa_tree_add_14_36_groupi_n_591 ();
drwire csa_tree_add_14_36_groupi_n_592 ();
drwire csa_tree_add_14_36_groupi_n_593 ();
drwire csa_tree_add_14_36_groupi_n_594 ();
drwire csa_tree_add_14_36_groupi_n_595 ();
drwire csa_tree_add_14_36_groupi_n_596 ();
drwire csa_tree_add_14_36_groupi_n_597 ();
drwire csa_tree_add_14_36_groupi_n_598 ();
drwire csa_tree_add_14_36_groupi_n_599 ();
drwire csa_tree_add_14_36_groupi_n_6 ();
drwire csa_tree_add_14_36_groupi_n_60 ();
drwire csa_tree_add_14_36_groupi_n_600 ();
drwire csa_tree_add_14_36_groupi_n_601 ();
drwire csa_tree_add_14_36_groupi_n_602 ();
drwire csa_tree_add_14_36_groupi_n_603 ();
drwire csa_tree_add_14_36_groupi_n_604 ();
drwire csa_tree_add_14_36_groupi_n_605 ();
drwire csa_tree_add_14_36_groupi_n_606 ();
drwire csa_tree_add_14_36_groupi_n_607 ();
drwire csa_tree_add_14_36_groupi_n_608 ();
drwire csa_tree_add_14_36_groupi_n_609 ();
drwire csa_tree_add_14_36_groupi_n_61 ();
drwire csa_tree_add_14_36_groupi_n_610 ();
drwire csa_tree_add_14_36_groupi_n_611 ();
drwire csa_tree_add_14_36_groupi_n_612 ();
drwire csa_tree_add_14_36_groupi_n_613 ();
drwire csa_tree_add_14_36_groupi_n_614 ();
drwire csa_tree_add_14_36_groupi_n_615 ();
drwire csa_tree_add_14_36_groupi_n_617 ();
drwire csa_tree_add_14_36_groupi_n_618 ();
drwire csa_tree_add_14_36_groupi_n_619 ();
drwire csa_tree_add_14_36_groupi_n_62 ();
drwire csa_tree_add_14_36_groupi_n_620 ();
drwire csa_tree_add_14_36_groupi_n_621 ();
drwire csa_tree_add_14_36_groupi_n_622 ();
drwire csa_tree_add_14_36_groupi_n_623 ();
drwire csa_tree_add_14_36_groupi_n_624 ();
drwire csa_tree_add_14_36_groupi_n_625 ();
drwire csa_tree_add_14_36_groupi_n_626 ();
drwire csa_tree_add_14_36_groupi_n_627 ();
drwire csa_tree_add_14_36_groupi_n_628 ();
drwire csa_tree_add_14_36_groupi_n_629 ();
drwire csa_tree_add_14_36_groupi_n_63 ();
drwire csa_tree_add_14_36_groupi_n_630 ();
drwire csa_tree_add_14_36_groupi_n_631 ();
drwire csa_tree_add_14_36_groupi_n_632 ();
drwire csa_tree_add_14_36_groupi_n_633 ();
drwire csa_tree_add_14_36_groupi_n_634 ();
drwire csa_tree_add_14_36_groupi_n_635 ();
drwire csa_tree_add_14_36_groupi_n_636 ();
drwire csa_tree_add_14_36_groupi_n_637 ();
drwire csa_tree_add_14_36_groupi_n_638 ();
drwire csa_tree_add_14_36_groupi_n_639 ();
drwire csa_tree_add_14_36_groupi_n_64 ();
drwire csa_tree_add_14_36_groupi_n_640 ();
drwire csa_tree_add_14_36_groupi_n_641 ();
drwire csa_tree_add_14_36_groupi_n_642 ();
drwire csa_tree_add_14_36_groupi_n_643 ();
drwire csa_tree_add_14_36_groupi_n_644 ();
drwire csa_tree_add_14_36_groupi_n_645 ();
drwire csa_tree_add_14_36_groupi_n_646 ();
drwire csa_tree_add_14_36_groupi_n_647 ();
drwire csa_tree_add_14_36_groupi_n_648 ();
drwire csa_tree_add_14_36_groupi_n_649 ();
drwire csa_tree_add_14_36_groupi_n_65 ();
drwire csa_tree_add_14_36_groupi_n_650 ();
drwire csa_tree_add_14_36_groupi_n_651 ();
drwire csa_tree_add_14_36_groupi_n_653 ();
drwire csa_tree_add_14_36_groupi_n_654 ();
drwire csa_tree_add_14_36_groupi_n_655 ();
drwire csa_tree_add_14_36_groupi_n_656 ();
drwire csa_tree_add_14_36_groupi_n_657 ();
drwire csa_tree_add_14_36_groupi_n_658 ();
drwire csa_tree_add_14_36_groupi_n_660 ();
drwire csa_tree_add_14_36_groupi_n_661 ();
drwire csa_tree_add_14_36_groupi_n_662 ();
drwire csa_tree_add_14_36_groupi_n_663 ();
drwire csa_tree_add_14_36_groupi_n_664 ();
drwire csa_tree_add_14_36_groupi_n_665 ();
drwire csa_tree_add_14_36_groupi_n_666 ();
drwire csa_tree_add_14_36_groupi_n_667 ();
drwire csa_tree_add_14_36_groupi_n_668 ();
drwire csa_tree_add_14_36_groupi_n_669 ();
drwire csa_tree_add_14_36_groupi_n_67 ();
drwire csa_tree_add_14_36_groupi_n_670 ();
drwire csa_tree_add_14_36_groupi_n_671 ();
drwire csa_tree_add_14_36_groupi_n_672 ();
drwire csa_tree_add_14_36_groupi_n_673 ();
drwire csa_tree_add_14_36_groupi_n_674 ();
drwire csa_tree_add_14_36_groupi_n_675 ();
drwire csa_tree_add_14_36_groupi_n_676 ();
drwire csa_tree_add_14_36_groupi_n_677 ();
drwire csa_tree_add_14_36_groupi_n_678 ();
drwire csa_tree_add_14_36_groupi_n_679 ();
drwire csa_tree_add_14_36_groupi_n_680 ();
drwire csa_tree_add_14_36_groupi_n_681 ();
drwire csa_tree_add_14_36_groupi_n_682 ();
drwire csa_tree_add_14_36_groupi_n_683 ();
drwire csa_tree_add_14_36_groupi_n_684 ();
drwire csa_tree_add_14_36_groupi_n_685 ();
drwire csa_tree_add_14_36_groupi_n_686 ();
drwire csa_tree_add_14_36_groupi_n_687 ();
drwire csa_tree_add_14_36_groupi_n_688 ();
drwire csa_tree_add_14_36_groupi_n_689 ();
drwire csa_tree_add_14_36_groupi_n_69 ();
drwire csa_tree_add_14_36_groupi_n_690 ();
drwire csa_tree_add_14_36_groupi_n_692 ();
drwire csa_tree_add_14_36_groupi_n_693 ();
drwire csa_tree_add_14_36_groupi_n_694 ();
drwire csa_tree_add_14_36_groupi_n_695 ();
drwire csa_tree_add_14_36_groupi_n_697 ();
drwire csa_tree_add_14_36_groupi_n_698 ();
drwire csa_tree_add_14_36_groupi_n_699 ();
drwire csa_tree_add_14_36_groupi_n_7 ();
drwire csa_tree_add_14_36_groupi_n_70 ();
drwire csa_tree_add_14_36_groupi_n_701 ();
drwire csa_tree_add_14_36_groupi_n_702 ();
drwire csa_tree_add_14_36_groupi_n_703 ();
drwire csa_tree_add_14_36_groupi_n_704 ();
drwire csa_tree_add_14_36_groupi_n_705 ();
drwire csa_tree_add_14_36_groupi_n_706 ();
drwire csa_tree_add_14_36_groupi_n_707 ();
drwire csa_tree_add_14_36_groupi_n_708 ();
drwire csa_tree_add_14_36_groupi_n_709 ();
drwire csa_tree_add_14_36_groupi_n_710 ();
drwire csa_tree_add_14_36_groupi_n_711 ();
drwire csa_tree_add_14_36_groupi_n_712 ();
drwire csa_tree_add_14_36_groupi_n_713 ();
drwire csa_tree_add_14_36_groupi_n_714 ();
drwire csa_tree_add_14_36_groupi_n_715 ();
drwire csa_tree_add_14_36_groupi_n_716 ();
drwire csa_tree_add_14_36_groupi_n_717 ();
drwire csa_tree_add_14_36_groupi_n_718 ();
drwire csa_tree_add_14_36_groupi_n_719 ();
drwire csa_tree_add_14_36_groupi_n_72 ();
drwire csa_tree_add_14_36_groupi_n_720 ();
drwire csa_tree_add_14_36_groupi_n_721 ();
drwire csa_tree_add_14_36_groupi_n_722 ();
drwire csa_tree_add_14_36_groupi_n_723 ();
drwire csa_tree_add_14_36_groupi_n_724 ();
drwire csa_tree_add_14_36_groupi_n_725 ();
drwire csa_tree_add_14_36_groupi_n_726 ();
drwire csa_tree_add_14_36_groupi_n_727 ();
drwire csa_tree_add_14_36_groupi_n_728 ();
drwire csa_tree_add_14_36_groupi_n_729 ();
drwire csa_tree_add_14_36_groupi_n_73 ();
drwire csa_tree_add_14_36_groupi_n_730 ();
drwire csa_tree_add_14_36_groupi_n_731 ();
drwire csa_tree_add_14_36_groupi_n_732 ();
drwire csa_tree_add_14_36_groupi_n_736 ();
drwire csa_tree_add_14_36_groupi_n_738 ();
drwire csa_tree_add_14_36_groupi_n_74 ();
drwire csa_tree_add_14_36_groupi_n_740 ();
drwire csa_tree_add_14_36_groupi_n_741 ();
drwire csa_tree_add_14_36_groupi_n_743 ();
drwire csa_tree_add_14_36_groupi_n_744 ();
drwire csa_tree_add_14_36_groupi_n_746 ();
drwire csa_tree_add_14_36_groupi_n_748 ();
drwire csa_tree_add_14_36_groupi_n_749 ();
drwire csa_tree_add_14_36_groupi_n_75 ();
drwire csa_tree_add_14_36_groupi_n_750 ();
drwire csa_tree_add_14_36_groupi_n_751 ();
drwire csa_tree_add_14_36_groupi_n_752 ();
drwire csa_tree_add_14_36_groupi_n_753 ();
drwire csa_tree_add_14_36_groupi_n_754 ();
drwire csa_tree_add_14_36_groupi_n_755 ();
drwire csa_tree_add_14_36_groupi_n_756 ();
drwire csa_tree_add_14_36_groupi_n_757 ();
drwire csa_tree_add_14_36_groupi_n_758 ();
drwire csa_tree_add_14_36_groupi_n_759 ();
drwire csa_tree_add_14_36_groupi_n_76 ();
drwire csa_tree_add_14_36_groupi_n_760 ();
drwire csa_tree_add_14_36_groupi_n_761 ();
drwire csa_tree_add_14_36_groupi_n_762 ();
drwire csa_tree_add_14_36_groupi_n_763 ();
drwire csa_tree_add_14_36_groupi_n_764 ();
drwire csa_tree_add_14_36_groupi_n_765 ();
drwire csa_tree_add_14_36_groupi_n_766 ();
drwire csa_tree_add_14_36_groupi_n_767 ();
drwire csa_tree_add_14_36_groupi_n_768 ();
drwire csa_tree_add_14_36_groupi_n_769 ();
drwire csa_tree_add_14_36_groupi_n_77 ();
drwire csa_tree_add_14_36_groupi_n_770 ();
drwire csa_tree_add_14_36_groupi_n_771 ();
drwire csa_tree_add_14_36_groupi_n_774 ();
drwire csa_tree_add_14_36_groupi_n_775 ();
drwire csa_tree_add_14_36_groupi_n_776 ();
drwire csa_tree_add_14_36_groupi_n_777 ();
drwire csa_tree_add_14_36_groupi_n_778 ();
drwire csa_tree_add_14_36_groupi_n_779 ();
drwire csa_tree_add_14_36_groupi_n_78 ();
drwire csa_tree_add_14_36_groupi_n_780 ();
drwire csa_tree_add_14_36_groupi_n_781 ();
drwire csa_tree_add_14_36_groupi_n_782 ();
drwire csa_tree_add_14_36_groupi_n_783 ();
drwire csa_tree_add_14_36_groupi_n_784 ();
drwire csa_tree_add_14_36_groupi_n_785 ();
drwire csa_tree_add_14_36_groupi_n_786 ();
drwire csa_tree_add_14_36_groupi_n_787 ();
drwire csa_tree_add_14_36_groupi_n_788 ();
drwire csa_tree_add_14_36_groupi_n_789 ();
drwire csa_tree_add_14_36_groupi_n_79 ();
drwire csa_tree_add_14_36_groupi_n_790 ();
drwire csa_tree_add_14_36_groupi_n_791 ();
drwire csa_tree_add_14_36_groupi_n_792 ();
drwire csa_tree_add_14_36_groupi_n_793 ();
drwire csa_tree_add_14_36_groupi_n_794 ();
drwire csa_tree_add_14_36_groupi_n_796 ();
drwire csa_tree_add_14_36_groupi_n_798 ();
drwire csa_tree_add_14_36_groupi_n_799 ();
drwire csa_tree_add_14_36_groupi_n_8 ();
drwire csa_tree_add_14_36_groupi_n_80 ();
drwire csa_tree_add_14_36_groupi_n_800 ();
drwire csa_tree_add_14_36_groupi_n_801 ();
drwire csa_tree_add_14_36_groupi_n_802 ();
drwire csa_tree_add_14_36_groupi_n_803 ();
drwire csa_tree_add_14_36_groupi_n_805 ();
drwire csa_tree_add_14_36_groupi_n_806 ();
drwire csa_tree_add_14_36_groupi_n_807 ();
drwire csa_tree_add_14_36_groupi_n_808 ();
drwire csa_tree_add_14_36_groupi_n_81 ();
drwire csa_tree_add_14_36_groupi_n_810 ();
drwire csa_tree_add_14_36_groupi_n_812 ();
drwire csa_tree_add_14_36_groupi_n_813 ();
drwire csa_tree_add_14_36_groupi_n_814 ();
drwire csa_tree_add_14_36_groupi_n_816 ();
drwire csa_tree_add_14_36_groupi_n_817 ();
drwire csa_tree_add_14_36_groupi_n_818 ();
drwire csa_tree_add_14_36_groupi_n_819 ();
drwire csa_tree_add_14_36_groupi_n_82 ();
drwire csa_tree_add_14_36_groupi_n_820 ();
drwire csa_tree_add_14_36_groupi_n_821 ();
drwire csa_tree_add_14_36_groupi_n_822 ();
drwire csa_tree_add_14_36_groupi_n_823 ();
drwire csa_tree_add_14_36_groupi_n_824 ();
drwire csa_tree_add_14_36_groupi_n_825 ();
drwire csa_tree_add_14_36_groupi_n_826 ();
drwire csa_tree_add_14_36_groupi_n_827 ();
drwire csa_tree_add_14_36_groupi_n_828 ();
drwire csa_tree_add_14_36_groupi_n_829 ();
drwire csa_tree_add_14_36_groupi_n_83 ();
drwire csa_tree_add_14_36_groupi_n_830 ();
drwire csa_tree_add_14_36_groupi_n_831 ();
drwire csa_tree_add_14_36_groupi_n_832 ();
drwire csa_tree_add_14_36_groupi_n_833 ();
drwire csa_tree_add_14_36_groupi_n_834 ();
drwire csa_tree_add_14_36_groupi_n_835 ();
drwire csa_tree_add_14_36_groupi_n_836 ();
drwire csa_tree_add_14_36_groupi_n_837 ();
drwire csa_tree_add_14_36_groupi_n_838 ();
drwire csa_tree_add_14_36_groupi_n_839 ();
drwire csa_tree_add_14_36_groupi_n_84 ();
drwire csa_tree_add_14_36_groupi_n_840 ();
drwire csa_tree_add_14_36_groupi_n_841 ();
drwire csa_tree_add_14_36_groupi_n_842 ();
drwire csa_tree_add_14_36_groupi_n_843 ();
drwire csa_tree_add_14_36_groupi_n_844 ();
drwire csa_tree_add_14_36_groupi_n_845 ();
drwire csa_tree_add_14_36_groupi_n_846 ();
drwire csa_tree_add_14_36_groupi_n_847 ();
drwire csa_tree_add_14_36_groupi_n_848 ();
drwire csa_tree_add_14_36_groupi_n_849 ();
drwire csa_tree_add_14_36_groupi_n_85 ();
drwire csa_tree_add_14_36_groupi_n_850 ();
drwire csa_tree_add_14_36_groupi_n_851 ();
drwire csa_tree_add_14_36_groupi_n_852 ();
drwire csa_tree_add_14_36_groupi_n_853 ();
drwire csa_tree_add_14_36_groupi_n_854 ();
drwire csa_tree_add_14_36_groupi_n_855 ();
drwire csa_tree_add_14_36_groupi_n_856 ();
drwire csa_tree_add_14_36_groupi_n_857 ();
drwire csa_tree_add_14_36_groupi_n_858 ();
drwire csa_tree_add_14_36_groupi_n_859 ();
drwire csa_tree_add_14_36_groupi_n_86 ();
drwire csa_tree_add_14_36_groupi_n_860 ();
drwire csa_tree_add_14_36_groupi_n_861 ();
drwire csa_tree_add_14_36_groupi_n_862 ();
drwire csa_tree_add_14_36_groupi_n_863 ();
drwire csa_tree_add_14_36_groupi_n_864 ();
drwire csa_tree_add_14_36_groupi_n_865 ();
drwire csa_tree_add_14_36_groupi_n_866 ();
drwire csa_tree_add_14_36_groupi_n_867 ();
drwire csa_tree_add_14_36_groupi_n_868 ();
drwire csa_tree_add_14_36_groupi_n_869 ();
drwire csa_tree_add_14_36_groupi_n_87 ();
drwire csa_tree_add_14_36_groupi_n_870 ();
drwire csa_tree_add_14_36_groupi_n_871 ();
drwire csa_tree_add_14_36_groupi_n_872 ();
drwire csa_tree_add_14_36_groupi_n_873 ();
drwire csa_tree_add_14_36_groupi_n_874 ();
drwire csa_tree_add_14_36_groupi_n_875 ();
drwire csa_tree_add_14_36_groupi_n_876 ();
drwire csa_tree_add_14_36_groupi_n_877 ();
drwire csa_tree_add_14_36_groupi_n_878 ();
drwire csa_tree_add_14_36_groupi_n_879 ();
drwire csa_tree_add_14_36_groupi_n_88 ();
drwire csa_tree_add_14_36_groupi_n_880 ();
drwire csa_tree_add_14_36_groupi_n_881 ();
drwire csa_tree_add_14_36_groupi_n_882 ();
drwire csa_tree_add_14_36_groupi_n_883 ();
drwire csa_tree_add_14_36_groupi_n_884 ();
drwire csa_tree_add_14_36_groupi_n_885 ();
drwire csa_tree_add_14_36_groupi_n_886 ();
drwire csa_tree_add_14_36_groupi_n_887 ();
drwire csa_tree_add_14_36_groupi_n_888 ();
drwire csa_tree_add_14_36_groupi_n_889 ();
drwire csa_tree_add_14_36_groupi_n_89 ();
drwire csa_tree_add_14_36_groupi_n_890 ();
drwire csa_tree_add_14_36_groupi_n_891 ();
drwire csa_tree_add_14_36_groupi_n_892 ();
drwire csa_tree_add_14_36_groupi_n_894 ();
drwire csa_tree_add_14_36_groupi_n_895 ();
drwire csa_tree_add_14_36_groupi_n_896 ();
drwire csa_tree_add_14_36_groupi_n_897 ();
drwire csa_tree_add_14_36_groupi_n_898 ();
drwire csa_tree_add_14_36_groupi_n_9 ();
drwire csa_tree_add_14_36_groupi_n_90 ();
drwire csa_tree_add_14_36_groupi_n_900 ();
drwire csa_tree_add_14_36_groupi_n_901 ();
drwire csa_tree_add_14_36_groupi_n_902 ();
drwire csa_tree_add_14_36_groupi_n_903 ();
drwire csa_tree_add_14_36_groupi_n_904 ();
drwire csa_tree_add_14_36_groupi_n_905 ();
drwire csa_tree_add_14_36_groupi_n_906 ();
drwire csa_tree_add_14_36_groupi_n_907 ();
drwire csa_tree_add_14_36_groupi_n_908 ();
drwire csa_tree_add_14_36_groupi_n_909 ();
drwire csa_tree_add_14_36_groupi_n_91 ();
drwire csa_tree_add_14_36_groupi_n_910 ();
drwire csa_tree_add_14_36_groupi_n_911 ();
drwire csa_tree_add_14_36_groupi_n_912 ();
drwire csa_tree_add_14_36_groupi_n_913 ();
drwire csa_tree_add_14_36_groupi_n_915 ();
drwire csa_tree_add_14_36_groupi_n_916 ();
drwire csa_tree_add_14_36_groupi_n_917 ();
drwire csa_tree_add_14_36_groupi_n_918 ();
drwire csa_tree_add_14_36_groupi_n_919 ();
drwire csa_tree_add_14_36_groupi_n_92 ();
drwire csa_tree_add_14_36_groupi_n_920 ();
drwire csa_tree_add_14_36_groupi_n_921 ();
drwire csa_tree_add_14_36_groupi_n_922 ();
drwire csa_tree_add_14_36_groupi_n_923 ();
drwire csa_tree_add_14_36_groupi_n_924 ();
drwire csa_tree_add_14_36_groupi_n_93 ();
drwire csa_tree_add_14_36_groupi_n_930 ();
drwire csa_tree_add_14_36_groupi_n_931 ();
drwire csa_tree_add_14_36_groupi_n_932 ();
drwire csa_tree_add_14_36_groupi_n_933 ();
drwire csa_tree_add_14_36_groupi_n_934 ();
drwire csa_tree_add_14_36_groupi_n_935 ();
drwire csa_tree_add_14_36_groupi_n_936 ();
drwire csa_tree_add_14_36_groupi_n_937 ();
drwire csa_tree_add_14_36_groupi_n_938 ();
drwire csa_tree_add_14_36_groupi_n_939 ();
drwire csa_tree_add_14_36_groupi_n_94 ();
drwire csa_tree_add_14_36_groupi_n_940 ();
drwire csa_tree_add_14_36_groupi_n_941 ();
drwire csa_tree_add_14_36_groupi_n_942 ();
drwire csa_tree_add_14_36_groupi_n_943 ();
drwire csa_tree_add_14_36_groupi_n_944 ();
drwire csa_tree_add_14_36_groupi_n_945 ();
drwire csa_tree_add_14_36_groupi_n_946 ();
drwire csa_tree_add_14_36_groupi_n_947 ();
drwire csa_tree_add_14_36_groupi_n_948 ();
drwire csa_tree_add_14_36_groupi_n_949 ();
drwire csa_tree_add_14_36_groupi_n_95 ();
drwire csa_tree_add_14_36_groupi_n_950 ();
drwire csa_tree_add_14_36_groupi_n_951 ();
drwire csa_tree_add_14_36_groupi_n_952 ();
drwire csa_tree_add_14_36_groupi_n_953 ();
drwire csa_tree_add_14_36_groupi_n_954 ();
drwire csa_tree_add_14_36_groupi_n_955 ();
drwire csa_tree_add_14_36_groupi_n_956 ();
drwire csa_tree_add_14_36_groupi_n_957 ();
drwire csa_tree_add_14_36_groupi_n_958 ();
drwire csa_tree_add_14_36_groupi_n_959 ();
drwire csa_tree_add_14_36_groupi_n_960 ();
drwire csa_tree_add_14_36_groupi_n_961 ();
drwire csa_tree_add_14_36_groupi_n_962 ();
drwire csa_tree_add_14_36_groupi_n_963 ();
drwire csa_tree_add_14_36_groupi_n_964 ();
drwire csa_tree_add_14_36_groupi_n_965 ();
drwire csa_tree_add_14_36_groupi_n_966 ();
drwire csa_tree_add_14_36_groupi_n_967 ();
drwire csa_tree_add_14_36_groupi_n_968 ();
drwire csa_tree_add_14_36_groupi_n_969 ();
drwire csa_tree_add_14_36_groupi_n_97 ();
drwire csa_tree_add_14_36_groupi_n_970 ();
drwire csa_tree_add_14_36_groupi_n_972 ();
drwire csa_tree_add_14_36_groupi_n_973 ();
drwire csa_tree_add_14_36_groupi_n_974 ();
drwire csa_tree_add_14_36_groupi_n_975 ();
drwire csa_tree_add_14_36_groupi_n_976 ();
drwire csa_tree_add_14_36_groupi_n_979 ();
drwire csa_tree_add_14_36_groupi_n_98 ();
drwire csa_tree_add_14_36_groupi_n_980 ();
drwire csa_tree_add_14_36_groupi_n_981 ();
drwire csa_tree_add_14_36_groupi_n_983 ();
drwire csa_tree_add_14_36_groupi_n_984 ();
drwire csa_tree_add_14_36_groupi_n_985 ();
drwire csa_tree_add_14_36_groupi_n_986 ();
drwire csa_tree_add_14_36_groupi_n_988 ();
drwire csa_tree_add_14_36_groupi_n_989 ();
drwire csa_tree_add_14_36_groupi_n_99 ();
drwire csa_tree_add_14_36_groupi_n_990 ();
drwire csa_tree_add_14_36_groupi_n_991 ();
drwire csa_tree_add_14_36_groupi_n_992 ();
drwire csa_tree_add_14_36_groupi_n_993 ();
drwire csa_tree_add_14_36_groupi_n_994 ();
drwire csa_tree_add_14_36_groupi_n_995 ();
drwire csa_tree_add_14_36_groupi_n_996 ();
drwire csa_tree_add_14_36_groupi_n_997 ();
drwire csa_tree_add_14_36_groupi_n_998 ();
drwire csa_tree_add_14_36_groupi_n_999 ();
drwire n_101 ();
drwire n_104 ();
drwire n_107 ();
drwire n_110 ();
drwire n_113 ();
drwire n_116 ();
drwire n_121 ();
drwire n_123 ();
drwire n_125 ();
drwire n_127 ();
drwire n_129 ();
drwire n_131 ();
drwire n_133 ();
drwire n_135 ();
drwire n_137 ();
drwire n_139 ();
drwire n_141 ();
drwire n_143 ();
drwire n_145 ();
drwire n_147 ();
drwire n_149 ();
drwire n_151 ();
drwire n_153 ();
drwire n_155 ();
drwire n_157 ();
drwire n_159 ();
drwire n_16 ();
drwire n_17 ();
drwire n_18 ();
drwire n_19 ();
drwire n_20 ();
drwire n_21 ();
drwire n_22 ();
drwire n_2424 ();
drwire n_2425 ();
drwire n_2426 ();
drwire n_2427 ();
drwire n_2428 ();
drwire n_2429 ();
drwire n_2430 ();
drwire n_2431 ();
drwire n_2432 ();
drwire n_2433 ();
drwire n_2434 ();
drwire n_2435 ();
drwire n_2436 ();
drwire n_2437 ();
drwire n_2438 ();
drwire n_2440 ();
drwire n_2445 ();
drwire n_2450 ();
drwire n_2451 ();
drwire n_2453 ();
drwire n_2455 ();
drwire n_2457 ();
drwire n_2458 ();
drwire n_2459 ();
drwire n_2460 ();
drwire n_2461 ();
drwire n_2462 ();
drwire n_2463 ();
drwire n_2464 ();
drwire n_2465 ();
drwire n_2466 ();
drwire n_2467 ();
drwire n_2468 ();
drwire n_2469 ();
drwire n_2470 ();
drwire n_2471 ();
drwire n_2472 ();
drwire n_2475 ();
drwire n_2476 ();
drwire n_2477 ();
drwire n_2478 ();
drwire n_2479 ();
drwire n_2480 ();
drwire n_2482 ();
drwire n_2483 ();
drwire n_2484 ();
drwire n_2485 ();
drwire n_2486 ();
drwire n_2487 ();
drwire n_2488 ();
drwire n_2489 ();
drwire n_2490 ();
drwire n_2491 ();
drwire n_2492 ();
drwire n_2503 ();
drwire n_2504 ();
drwire n_2505 ();
drwire n_2506 ();
drwire n_2507 ();
drwire n_2508 ();
drwire n_2509 ();
drwire n_2510 ();
drwire n_2511 ();
drwire n_2513 ();
drwire n_2514 ();
drwire n_2515 ();
drwire n_2516 ();
drwire n_2517 ();
drwire n_2518 ();
drwire n_2519 ();
drwire n_2520 ();
drwire n_2521 ();
drwire n_2522 ();
drwire n_2523 ();
drwire n_2524 ();
drwire n_2525 ();
drwire n_2526 ();
drwire n_2527 ();
drwire n_2528 ();
drwire n_2529 ();
drwire n_2537 ();
drwire n_2542 ();
drwire n_2543 ();
drwire n_2544 ();
drwire n_2546 ();
drwire n_2547 ();
drwire n_2548 ();
drwire n_2549 ();
drwire n_2550 ();
drwire n_2551 ();
drwire n_2553 ();
drwire n_2554 ();
drwire n_2556 ();
drwire n_2558 ();
drwire n_2559 ();
drwire n_2561 ();
drwire n_2564 ();
drwire n_2565 ();
drwire n_2566 ();
drwire n_2567 ();
drwire n_2568 ();
drwire n_2569 ();
drwire n_2570 ();
drwire n_2574 ();
drwire n_2575 ();
drwire n_2576 ();
drwire n_2577 ();
drwire n_2582 ();
drwire n_2583 ();
drwire n_2585 ();
drwire n_2586 ();
drwire n_2605 ();
drwire n_2606 ();
drwire n_2607 ();
drwire n_2609 ();
drwire n_2611 ();
drwire n_2612 ();
drwire n_2614 ();
drwire n_2616 ();
drwire n_2617 ();
drwire n_2618 ();
drwire n_2620 ();
drwire n_2621 ();
drwire n_2622 ();
drwire n_2623 ();
drwire n_2624 ();
drwire n_2631 ();
drwire n_2632 ();
drwire n_2633 ();
drwire n_2634 ();
drwire n_2635 ();
drwire n_2637 ();
drwire n_2638 ();
drwire n_2639 ();
drwire n_2640 ();
drwire n_2641 ();
drwire n_2642 ();
drwire n_2643 ();
drwire n_2644 ();
drwire n_2645 ();
drwire n_2646 ();
drwire n_2654 ();
drwire n_2655 ();
drwire n_2656 ();
drwire n_2657 ();
drwire n_2658 ();
drwire n_2659 ();
drwire n_2673 ();
drwire n_2674 ();
drwire n_2675 ();
drwire n_2676 ();
drwire n_2677 ();
drwire n_2678 ();
drwire n_2681 ();
drwire n_2682 ();
drwire n_2683 ();
drwire n_2684 ();
drwire n_2685 ();
drwire n_2687 ();
drwire n_2688 ();
drwire n_2689 ();
drwire n_2690 ();
drwire n_2693 ();
drwire n_2695 ();
drwire n_2696 ();
drwire n_2697 ();
drwire n_2698 ();
drwire n_2751 ();
drwire n_2752 ();
drwire n_2753 ();
drwire n_2754 ();
drwire n_2755 ();
drwire n_2756 ();
drwire n_2757 ();
drwire n_2758 ();
drwire n_2759 ();
drwire n_2760 ();
drwire n_2761 ();
drwire n_2762 ();
drwire n_2763 ();
drwire n_2764 ();
drwire n_2765 ();
drwire n_2766 ();
drwire n_2767 ();
drwire n_2768 ();
drwire n_2769 ();
drwire n_2770 ();
drwire n_2771 ();
drwire n_2772 ();
drwire n_2774 ();
drwire n_2775 ();
drwire n_2776 ();
drwire n_2777 ();
drwire n_2778 ();
drwire n_2779 ();
drwire n_2780 ();
drwire n_2781 ();
drwire n_75 ();
drwire n_76 ();
drwire n_77 ();
drwire n_78 ();
drwire n_79 ();
drwire n_80 ();
drwire n_81 ();
drwire n_82 ();
drwire n_83 ();
drwire n_84 ();
drwire n_85 ();
drwire n_86 ();
drwire n_89 ();
drwire n_92 ();
drwire n_95 ();
drwire n_98 ();
drwire result_0__0_ ();
drwire result_0__10_ ();
drwire result_0__11_ ();
drwire result_0__12_ ();
drwire result_0__13_ ();
drwire result_0__14_ ();
drwire result_0__15_ ();
drwire result_0__16_ ();
drwire result_0__17_ ();
drwire result_0__18_ ();
drwire result_0__19_ ();
drwire result_0__1_ ();
drwire result_0__20_ ();
drwire result_0__21_ ();
drwire result_0__22_ ();
drwire result_0__23_ ();
drwire result_0__24_ ();
drwire result_0__25_ ();
drwire result_0__26_ ();
drwire result_0__27_ ();
drwire result_0__28_ ();
drwire result_0__29_ ();
drwire result_0__2_ ();
drwire result_0__30_ ();
drwire result_0__31_ ();
drwire result_0__3_ ();
drwire result_0__4_ ();
drwire result_0__5_ ();
drwire result_0__6_ ();
drwire result_0__7_ ();
drwire result_0__8_ ();
drwire result_0__9_ ();
drwire a_0 ();
drwire a_1 ();
drwire a_2 ();
drwire a_3 ();
drwire a_4 ();
drwire a_5 ();
drwire a_6 ();
drwire a_7 ();
drwire a_8 ();
drwire a_9 ();
drwire a_10 ();
drwire a_11 ();
drwire a_12 ();
drwire a_13 ();
drwire a_14 ();
drwire a_15 ();
drwire b_0 ();
drwire b_1 ();
drwire b_2 ();
drwire b_3 ();
drwire b_4 ();
drwire b_5 ();
drwire b_6 ();
drwire b_7 ();
drwire b_8 ();
drwire b_9 ();
drwire b_10 ();
drwire b_11 ();
drwire b_12 ();
drwire b_13 ();
drwire b_14 ();
drwire b_15 ();
drwire out_0 ();
drwire out_1 ();
drwire out_2 ();
drwire out_3 ();
drwire out_4 ();
drwire out_5 ();
drwire out_6 ();
drwire out_7 ();
drwire out_8 ();
drwire out_9 ();
drwire out_10 ();
drwire out_11 ();
drwire out_12 ();
drwire out_13 ();
drwire out_14 ();
drwire out_15 ();
drwire out_16 ();
drwire out_17 ();
drwire out_18 ();
drwire out_19 ();
drwire out_20 ();
drwire out_21 ();
drwire out_22 ();
drwire out_23 ();
drwire out_24 ();
drwire out_25 ();
drwire out_26 ();
drwire out_27 ();
drwire out_28 ();
drwire out_29 ();
drwire out_30 ();
drwire out_31 ();
input  [15:0] a_t, a_f;
output [15:0] a_ack;
drinput ia_0 (.t(a_t[0]), .f(a_f[0]), .ack(a_ack[0]), .drw(a_0));
drinput ia_1 (.t(a_t[1]), .f(a_f[1]), .ack(a_ack[1]), .drw(a_1));
drinput ia_2 (.t(a_t[2]), .f(a_f[2]), .ack(a_ack[2]), .drw(a_2));
drinput ia_3 (.t(a_t[3]), .f(a_f[3]), .ack(a_ack[3]), .drw(a_3));
drinput ia_4 (.t(a_t[4]), .f(a_f[4]), .ack(a_ack[4]), .drw(a_4));
drinput ia_5 (.t(a_t[5]), .f(a_f[5]), .ack(a_ack[5]), .drw(a_5));
drinput ia_6 (.t(a_t[6]), .f(a_f[6]), .ack(a_ack[6]), .drw(a_6));
drinput ia_7 (.t(a_t[7]), .f(a_f[7]), .ack(a_ack[7]), .drw(a_7));
drinput ia_8 (.t(a_t[8]), .f(a_f[8]), .ack(a_ack[8]), .drw(a_8));
drinput ia_9 (.t(a_t[9]), .f(a_f[9]), .ack(a_ack[9]), .drw(a_9));
drinput ia_10 (.t(a_t[10]), .f(a_f[10]), .ack(a_ack[10]), .drw(a_10));
drinput ia_11 (.t(a_t[11]), .f(a_f[11]), .ack(a_ack[11]), .drw(a_11));
drinput ia_12 (.t(a_t[12]), .f(a_f[12]), .ack(a_ack[12]), .drw(a_12));
drinput ia_13 (.t(a_t[13]), .f(a_f[13]), .ack(a_ack[13]), .drw(a_13));
drinput ia_14 (.t(a_t[14]), .f(a_f[14]), .ack(a_ack[14]), .drw(a_14));
drinput ia_15 (.t(a_t[15]), .f(a_f[15]), .ack(a_ack[15]), .drw(a_15));
input  [15:0] b_t, b_f;
output [15:0] b_ack;
drinput ib_0 (.t(b_t[0]), .f(b_f[0]), .ack(b_ack[0]), .drw(b_0));
drinput ib_1 (.t(b_t[1]), .f(b_f[1]), .ack(b_ack[1]), .drw(b_1));
drinput ib_2 (.t(b_t[2]), .f(b_f[2]), .ack(b_ack[2]), .drw(b_2));
drinput ib_3 (.t(b_t[3]), .f(b_f[3]), .ack(b_ack[3]), .drw(b_3));
drinput ib_4 (.t(b_t[4]), .f(b_f[4]), .ack(b_ack[4]), .drw(b_4));
drinput ib_5 (.t(b_t[5]), .f(b_f[5]), .ack(b_ack[5]), .drw(b_5));
drinput ib_6 (.t(b_t[6]), .f(b_f[6]), .ack(b_ack[6]), .drw(b_6));
drinput ib_7 (.t(b_t[7]), .f(b_f[7]), .ack(b_ack[7]), .drw(b_7));
drinput ib_8 (.t(b_t[8]), .f(b_f[8]), .ack(b_ack[8]), .drw(b_8));
drinput ib_9 (.t(b_t[9]), .f(b_f[9]), .ack(b_ack[9]), .drw(b_9));
drinput ib_10 (.t(b_t[10]), .f(b_f[10]), .ack(b_ack[10]), .drw(b_10));
drinput ib_11 (.t(b_t[11]), .f(b_f[11]), .ack(b_ack[11]), .drw(b_11));
drinput ib_12 (.t(b_t[12]), .f(b_f[12]), .ack(b_ack[12]), .drw(b_12));
drinput ib_13 (.t(b_t[13]), .f(b_f[13]), .ack(b_ack[13]), .drw(b_13));
drinput ib_14 (.t(b_t[14]), .f(b_f[14]), .ack(b_ack[14]), .drw(b_14));
drinput ib_15 (.t(b_t[15]), .f(b_f[15]), .ack(b_ack[15]), .drw(b_15));
output [31:0] out_t, out_f;
input  [31:0] out_ack;
droutput iout_0 (.t(out_t[0]), .f(out_f[0]), .ack(out_ack[0]), .drw(out_0));
droutput iout_1 (.t(out_t[1]), .f(out_f[1]), .ack(out_ack[1]), .drw(out_1));
droutput iout_2 (.t(out_t[2]), .f(out_f[2]), .ack(out_ack[2]), .drw(out_2));
droutput iout_3 (.t(out_t[3]), .f(out_f[3]), .ack(out_ack[3]), .drw(out_3));
droutput iout_4 (.t(out_t[4]), .f(out_f[4]), .ack(out_ack[4]), .drw(out_4));
droutput iout_5 (.t(out_t[5]), .f(out_f[5]), .ack(out_ack[5]), .drw(out_5));
droutput iout_6 (.t(out_t[6]), .f(out_f[6]), .ack(out_ack[6]), .drw(out_6));
droutput iout_7 (.t(out_t[7]), .f(out_f[7]), .ack(out_ack[7]), .drw(out_7));
droutput iout_8 (.t(out_t[8]), .f(out_f[8]), .ack(out_ack[8]), .drw(out_8));
droutput iout_9 (.t(out_t[9]), .f(out_f[9]), .ack(out_ack[9]), .drw(out_9));
droutput iout_10 (.t(out_t[10]), .f(out_f[10]), .ack(out_ack[10]), .drw(out_10));
droutput iout_11 (.t(out_t[11]), .f(out_f[11]), .ack(out_ack[11]), .drw(out_11));
droutput iout_12 (.t(out_t[12]), .f(out_f[12]), .ack(out_ack[12]), .drw(out_12));
droutput iout_13 (.t(out_t[13]), .f(out_f[13]), .ack(out_ack[13]), .drw(out_13));
droutput iout_14 (.t(out_t[14]), .f(out_f[14]), .ack(out_ack[14]), .drw(out_14));
droutput iout_15 (.t(out_t[15]), .f(out_f[15]), .ack(out_ack[15]), .drw(out_15));
droutput iout_16 (.t(out_t[16]), .f(out_f[16]), .ack(out_ack[16]), .drw(out_16));
droutput iout_17 (.t(out_t[17]), .f(out_f[17]), .ack(out_ack[17]), .drw(out_17));
droutput iout_18 (.t(out_t[18]), .f(out_f[18]), .ack(out_ack[18]), .drw(out_18));
droutput iout_19 (.t(out_t[19]), .f(out_f[19]), .ack(out_ack[19]), .drw(out_19));
droutput iout_20 (.t(out_t[20]), .f(out_f[20]), .ack(out_ack[20]), .drw(out_20));
droutput iout_21 (.t(out_t[21]), .f(out_f[21]), .ack(out_ack[21]), .drw(out_21));
droutput iout_22 (.t(out_t[22]), .f(out_f[22]), .ack(out_ack[22]), .drw(out_22));
droutput iout_23 (.t(out_t[23]), .f(out_f[23]), .ack(out_ack[23]), .drw(out_23));
droutput iout_24 (.t(out_t[24]), .f(out_f[24]), .ack(out_ack[24]), .drw(out_24));
droutput iout_25 (.t(out_t[25]), .f(out_f[25]), .ack(out_ack[25]), .drw(out_25));
droutput iout_26 (.t(out_t[26]), .f(out_f[26]), .ack(out_ack[26]), .drw(out_26));
droutput iout_27 (.t(out_t[27]), .f(out_f[27]), .ack(out_ack[27]), .drw(out_27));
droutput iout_28 (.t(out_t[28]), .f(out_f[28]), .ack(out_ack[28]), .drw(out_28));
droutput iout_29 (.t(out_t[29]), .f(out_f[29]), .ack(out_ack[29]), .drw(out_29));
droutput iout_30 (.t(out_t[30]), .f(out_f[30]), .ack(out_ack[30]), .drw(out_30));
droutput iout_31 (.t(out_t[31]), .f(out_f[31]), .ack(out_ack[31]), .drw(out_31));
dffr retime_s7_1_reg (.rb(reset), .ck(clk), .d(n_22), .q(n_75));
dffr retime_s4_1_reg (.rb(reset), .ck(clk), .d(n_21), .q(n_76));
dff retime_s3_6_reg (.reset(reset), .ck(clk), .d(n_20), .q(n_101));
dff retime_s3_8_reg (.reset(reset), .ck(clk), .d(n_18), .q(n_95));
dff retime_s4_2_reg (.reset(reset), .ck(clk), .d(n_21), .q(out_10));
dff retime_s7_2_reg (.reset(reset), .ck(clk), .d(n_22), .q(out_12));
dff retime_s3_7_reg (.reset(reset), .ck(clk), .d(n_19), .q(n_98));
dff retime_s3_9_reg (.reset(reset), .ck(clk), .d(n_17), .q(n_92));
dff retime_s3_10_reg (.reset(reset), .ck(clk), .d(n_16), .q(n_89));
dff retime_s4_9_reg (.reset(reset), .ck(clk), .d(n_101), .q(out_4));
dffr acc_reg_17_ (.rb(reset), .ck(clk), .d(result_0__17_), .q(n_153));
dffr acc_reg_18_ (.rb(reset), .ck(clk), .d(result_0__18_), .q(n_125));
dffr acc_reg_22_ (.rb(reset), .ck(clk), .d(result_0__22_), .q(n_149));
dffr acc_reg_24_ (.rb(reset), .ck(clk), .d(result_0__24_), .q(n_147));
dffr acc_reg_25_ (.rb(reset), .ck(clk), .d(result_0__25_), .q(n_133));
dffr acc_reg_13_ (.rb(reset), .ck(clk), .d(result_0__13_), .q(n_157));
dffr acc_reg_31_ (.rb(reset), .ck(clk), .d(result_0__31_), .q(n_143));
dffr acc_reg_27_ (.rb(reset), .ck(clk), .d(result_0__27_), .q(n_141));
dff retime_s4_4_reg (.reset(reset), .ck(clk), .d(n_116), .q(out_9));
dff retime_s4_6_reg (.reset(reset), .ck(clk), .d(n_113), .q(out_8));
dff retime_s4_8_reg (.reset(reset), .ck(clk), .d(n_110), .q(out_5));
dffr acc_reg_16_ (.rb(reset), .ck(clk), .d(result_0__16_), .q(n_123));
dff retime_s4_13_reg (.reset(reset), .ck(clk), .d(n_95), .q(out_2));
dff retime_s4_11_reg (.reset(reset), .ck(clk), .d(n_98), .q(out_3));
dff retime_s4_15_reg (.reset(reset), .ck(clk), .d(n_92), .q(out_1));
dff retime_s4_17_reg (.reset(reset), .ck(clk), .d(n_89), .q(out_0));
dff retime_s7_6_reg (.reset(reset), .ck(clk), .d(n_104), .q(out_6));
dff retime_s7_4_reg (.reset(reset), .ck(clk), .d(n_107), .q(out_7));
dff retime_s2_7_reg (.reset(reset), .ck(clk), .d(result_0__3_), .q(n_19));
dff retime_s6_2_reg (.reset(reset), .ck(clk), .d(result_0__12_), .q(n_22));
dff retime_s6_4_reg (.reset(reset), .ck(clk), .d(result_0__7_), .q(n_107));
dff retime_s6_5_reg (.reset(reset), .ck(clk), .d(result_0__6_), .q(n_104));
dff retime_s3_2_reg (.reset(reset), .ck(clk), .d(result_0__10_), .q(n_21));
dff retime_s3_5_reg (.reset(reset), .ck(clk), .d(result_0__5_), .q(n_110));
dff out_reg_24_ (.reset(reset), .ck(clk), .d(result_0__24_), .q(out_24));
dff out_reg_13_ (.reset(reset), .ck(clk), .d(result_0__13_), .q(out_13));
dff out_reg_14_ (.reset(reset), .ck(clk), .d(result_0__14_), .q(out_14));
dff out_reg_15_ (.reset(reset), .ck(clk), .d(result_0__15_), .q(out_15));
dff out_reg_25_ (.reset(reset), .ck(clk), .d(result_0__25_), .q(out_25));
dff out_reg_16_ (.reset(reset), .ck(clk), .d(result_0__16_), .q(out_16));
dff out_reg_17_ (.reset(reset), .ck(clk), .d(result_0__17_), .q(out_17));
dff out_reg_18_ (.reset(reset), .ck(clk), .d(result_0__18_), .q(out_18));
dff out_reg_19_ (.reset(reset), .ck(clk), .d(result_0__19_), .q(out_19));
dff out_reg_20_ (.reset(reset), .ck(clk), .d(result_0__20_), .q(out_20));
dff out_reg_21_ (.reset(reset), .ck(clk), .d(result_0__21_), .q(out_21));
dff out_reg_22_ (.reset(reset), .ck(clk), .d(result_0__22_), .q(out_22));
dff out_reg_23_ (.reset(reset), .ck(clk), .d(result_0__23_), .q(out_23));
dff out_reg_11_ (.reset(reset), .ck(clk), .d(result_0__11_), .q(out_11));
dff out_reg_27_ (.reset(reset), .ck(clk), .d(result_0__27_), .q(out_27));
dff out_reg_28_ (.reset(reset), .ck(clk), .d(result_0__28_), .q(out_28));
dff out_reg_29_ (.reset(reset), .ck(clk), .d(result_0__29_), .q(out_29));
dff out_reg_30_ (.reset(reset), .ck(clk), .d(result_0__30_), .q(out_30));
dff out_reg_31_ (.reset(reset), .ck(clk), .d(result_0__31_), .q(out_31));
dff retime_s2_6_reg (.reset(reset), .ck(clk), .d(result_0__4_), .q(n_20));
dff out_reg_26_ (.reset(reset), .ck(clk), .d(result_0__26_), .q(out_26));
dff retime_s2_11_reg (.reset(reset), .ck(clk), .d(result_0__1_), .q(n_17));
dff retime_s2_13_reg (.reset(reset), .ck(clk), .d(result_0__0_), .q(n_16));
dff retime_s2_8_reg (.reset(reset), .ck(clk), .d(result_0__2_), .q(n_18));
dff retime_s3_3_reg (.reset(reset), .ck(clk), .d(result_0__9_), .q(n_116));
dff retime_s3_4_reg (.reset(reset), .ck(clk), .d(result_0__8_), .q(n_113));
dffr acc_reg_11_ (.rb(reset), .ck(clk), .d(result_0__11_), .q(n_159));
dffr acc_reg_14_ (.rb(reset), .ck(clk), .d(result_0__14_), .q(n_121));
dffr retime_s4_18_reg (.rb(reset), .ck(clk), .d(n_89), .q(n_86));
dffr retime_s7_3_reg (.rb(reset), .ck(clk), .d(n_107), .q(n_79));
dffr retime_s4_16_reg (.rb(reset), .ck(clk), .d(n_92), .q(n_85));
dffr retime_s7_5_reg (.rb(reset), .ck(clk), .d(n_104), .q(n_80));
dffr acc_reg_15_ (.rb(reset), .ck(clk), .d(result_0__15_), .q(n_155));
dffr acc_reg_19_ (.rb(reset), .ck(clk), .d(result_0__19_), .q(n_151));
dffr retime_s4_7_reg (.rb(reset), .ck(clk), .d(n_110), .q(n_81));
dffr acc_reg_20_ (.rb(reset), .ck(clk), .d(result_0__20_), .q(n_127));
dffr acc_reg_30_ (.rb(reset), .ck(clk), .d(result_0__30_), .q(n_135));
dffr acc_reg_23_ (.rb(reset), .ck(clk), .d(result_0__23_), .q(n_131));
dffr acc_reg_26_ (.rb(reset), .ck(clk), .d(result_0__26_), .q(n_139));
dffr acc_reg_28_ (.rb(reset), .ck(clk), .d(result_0__28_), .q(n_145));
dffr acc_reg_29_ (.rb(reset), .ck(clk), .d(result_0__29_), .q(n_137));
dffr acc_reg_21_ (.rb(reset), .ck(clk), .d(result_0__21_), .q(n_129));
dffr retime_s4_3_reg (.rb(reset), .ck(clk), .d(n_116), .q(n_77));
dffr retime_s4_5_reg (.rb(reset), .ck(clk), .d(n_113), .q(n_78));
dffr retime_s4_10_reg (.rb(reset), .ck(clk), .d(n_101), .q(n_82));
dffr retime_s4_12_reg (.rb(reset), .ck(clk), .d(n_98), .q(n_83));
dffr retime_s4_14_reg (.rb(reset), .ck(clk), .d(n_95), .q(n_84));
dff csa_tree_add_14_36_groupi_retime_s1_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_323), .q(csa_tree_add_14_36_groupi_n_2260));
dff csa_tree_add_14_36_groupi_retime_s1_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_89), .q(csa_tree_add_14_36_groupi_n_2304));
dff csa_tree_add_14_36_groupi_retime_s1_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_331), .q(csa_tree_add_14_36_groupi_n_2167));
dff csa_tree_add_14_36_groupi_retime_s1_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_94), .q(csa_tree_add_14_36_groupi_n_2158));
dff csa_tree_add_14_36_groupi_retime_s1_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_332), .q(csa_tree_add_14_36_groupi_n_2157));
dff csa_tree_add_14_36_groupi_retime_s1_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_329), .q(csa_tree_add_14_36_groupi_n_2156));
dff csa_tree_add_14_36_groupi_retime_s1_7_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_99), .q(csa_tree_add_14_36_groupi_n_2155));
dff csa_tree_add_14_36_groupi_retime_s1_8_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_333), .q(csa_tree_add_14_36_groupi_n_2154));
dff csa_tree_add_14_36_groupi_retime_s1_9_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_322), .q(csa_tree_add_14_36_groupi_n_2153));
dff csa_tree_add_14_36_groupi_retime_s1_10_reg (.reset(reset), .ck(clk), .d(n_2529), .q(csa_tree_add_14_36_groupi_n_2152));
dff csa_tree_add_14_36_groupi_retime_s1_11_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1166), .q(csa_tree_add_14_36_groupi_n_2151));
dff csa_tree_add_14_36_groupi_retime_s1_12_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_687), .q(csa_tree_add_14_36_groupi_n_2302));
dff csa_tree_add_14_36_groupi_retime_s1_13_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1110), .q(csa_tree_add_14_36_groupi_n_2150));
dff csa_tree_add_14_36_groupi_retime_s1_14_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_759), .q(csa_tree_add_14_36_groupi_n_2149));
dff csa_tree_add_14_36_groupi_retime_s1_15_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1152), .q(csa_tree_add_14_36_groupi_n_2148));
dff csa_tree_add_14_36_groupi_retime_s1_16_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1108), .q(csa_tree_add_14_36_groupi_n_2147));
dff csa_tree_add_14_36_groupi_retime_s1_17_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1169), .q(csa_tree_add_14_36_groupi_n_2146));
dff csa_tree_add_14_36_groupi_retime_s1_18_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1096), .q(csa_tree_add_14_36_groupi_n_2145));
dff csa_tree_add_14_36_groupi_retime_s1_19_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_665), .q(csa_tree_add_14_36_groupi_n_2144));
dff csa_tree_add_14_36_groupi_retime_s1_20_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_632), .q(csa_tree_add_14_36_groupi_n_2143));
dff csa_tree_add_14_36_groupi_retime_s1_21_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1488), .q(csa_tree_add_14_36_groupi_n_2142));
dff csa_tree_add_14_36_groupi_retime_s1_22_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_695), .q(csa_tree_add_14_36_groupi_n_2140));
dff csa_tree_add_14_36_groupi_retime_s1_23_reg (.reset(reset), .ck(clk), .d(n_2771), .q(csa_tree_add_14_36_groupi_n_2139));
dff csa_tree_add_14_36_groupi_retime_s1_24_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_672), .q(csa_tree_add_14_36_groupi_n_2137));
dff csa_tree_add_14_36_groupi_retime_s1_25_reg (.reset(reset), .ck(clk), .d(n_2618), .q(csa_tree_add_14_36_groupi_n_2136));
dff csa_tree_add_14_36_groupi_retime_s1_26_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_615), .q(csa_tree_add_14_36_groupi_n_2135));
dff csa_tree_add_14_36_groupi_retime_s1_27_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_698), .q(csa_tree_add_14_36_groupi_n_2134));
dff csa_tree_add_14_36_groupi_retime_s1_28_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1068), .q(csa_tree_add_14_36_groupi_n_2133));
dff csa_tree_add_14_36_groupi_retime_s1_29_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_932), .q(csa_tree_add_14_36_groupi_n_2132));
dff csa_tree_add_14_36_groupi_retime_s1_30_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_951), .q(csa_tree_add_14_36_groupi_n_2131));
dff csa_tree_add_14_36_groupi_retime_s1_31_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1490), .q(csa_tree_add_14_36_groupi_n_2130));
dff csa_tree_add_14_36_groupi_retime_s1_32_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1239), .q(csa_tree_add_14_36_groupi_n_2129));
dff csa_tree_add_14_36_groupi_retime_s1_33_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_694), .q(csa_tree_add_14_36_groupi_n_2128));
dff csa_tree_add_14_36_groupi_retime_s1_34_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1350), .q(csa_tree_add_14_36_groupi_n_2127));
dff csa_tree_add_14_36_groupi_retime_s1_35_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1114), .q(csa_tree_add_14_36_groupi_n_2126));
dff csa_tree_add_14_36_groupi_retime_s1_36_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_671), .q(csa_tree_add_14_36_groupi_n_2125));
dff csa_tree_add_14_36_groupi_retime_s1_37_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_501), .q(csa_tree_add_14_36_groupi_n_2124));
dff csa_tree_add_14_36_groupi_retime_s1_38_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_490), .q(csa_tree_add_14_36_groupi_n_2123));
dff csa_tree_add_14_36_groupi_retime_s1_39_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1116), .q(csa_tree_add_14_36_groupi_n_2301));
dff csa_tree_add_14_36_groupi_retime_s1_40_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1099), .q(csa_tree_add_14_36_groupi_n_2122));
dff csa_tree_add_14_36_groupi_retime_s1_41_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1246), .q(csa_tree_add_14_36_groupi_n_2121));
dff csa_tree_add_14_36_groupi_retime_s1_42_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1288), .q(csa_tree_add_14_36_groupi_n_2120));
dff csa_tree_add_14_36_groupi_retime_s1_43_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1164), .q(csa_tree_add_14_36_groupi_n_2119));
dff csa_tree_add_14_36_groupi_retime_s1_44_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1168), .q(csa_tree_add_14_36_groupi_n_2118));
dff csa_tree_add_14_36_groupi_retime_s1_45_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1151), .q(csa_tree_add_14_36_groupi_n_2117));
dff csa_tree_add_14_36_groupi_retime_s1_46_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_670), .q(csa_tree_add_14_36_groupi_n_2116));
dff csa_tree_add_14_36_groupi_retime_s1_47_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_526), .q(csa_tree_add_14_36_groupi_n_2115));
dff csa_tree_add_14_36_groupi_retime_s1_48_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1095), .q(csa_tree_add_14_36_groupi_n_2114));
dff csa_tree_add_14_36_groupi_retime_s1_49_reg (.reset(reset), .ck(clk), .d(n_2524), .q(csa_tree_add_14_36_groupi_n_2113));
dff csa_tree_add_14_36_groupi_retime_s1_50_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1074), .q(csa_tree_add_14_36_groupi_n_2112));
dff csa_tree_add_14_36_groupi_retime_s1_51_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1105), .q(csa_tree_add_14_36_groupi_n_2111));
dff csa_tree_add_14_36_groupi_retime_s1_52_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_758), .q(csa_tree_add_14_36_groupi_n_2110));
dff csa_tree_add_14_36_groupi_retime_s1_53_reg (.reset(reset), .ck(clk), .d(n_2519), .q(csa_tree_add_14_36_groupi_n_2300));
dff csa_tree_add_14_36_groupi_retime_s1_54_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1170), .q(csa_tree_add_14_36_groupi_n_2109));
dff csa_tree_add_14_36_groupi_retime_s1_55_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1098), .q(csa_tree_add_14_36_groupi_n_2108));
dff csa_tree_add_14_36_groupi_retime_s1_56_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1123), .q(csa_tree_add_14_36_groupi_n_2107));
dff csa_tree_add_14_36_groupi_retime_s1_57_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_528), .q(csa_tree_add_14_36_groupi_n_2106));
dff csa_tree_add_14_36_groupi_retime_s1_58_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_760), .q(csa_tree_add_14_36_groupi_n_2105));
dff csa_tree_add_14_36_groupi_retime_s1_59_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1172), .q(csa_tree_add_14_36_groupi_n_2104));
dff csa_tree_add_14_36_groupi_retime_s1_60_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_761), .q(csa_tree_add_14_36_groupi_n_2103));
dff csa_tree_add_14_36_groupi_retime_s1_61_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_762), .q(csa_tree_add_14_36_groupi_n_2102));
dff csa_tree_add_14_36_groupi_retime_s1_62_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1107), .q(csa_tree_add_14_36_groupi_n_2101));
dff csa_tree_add_14_36_groupi_retime_s1_63_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1171), .q(csa_tree_add_14_36_groupi_n_2299));
dff csa_tree_add_14_36_groupi_retime_s1_64_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1100), .q(csa_tree_add_14_36_groupi_n_2100));
dff csa_tree_add_14_36_groupi_retime_s1_65_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1162), .q(csa_tree_add_14_36_groupi_n_2099));
dff csa_tree_add_14_36_groupi_retime_s1_66_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1241), .q(csa_tree_add_14_36_groupi_n_2098));
dff csa_tree_add_14_36_groupi_retime_s1_67_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_689), .q(csa_tree_add_14_36_groupi_n_2096));
dff csa_tree_add_14_36_groupi_retime_s1_68_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1153), .q(csa_tree_add_14_36_groupi_n_2095));
dff csa_tree_add_14_36_groupi_retime_s1_69_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_664), .q(csa_tree_add_14_36_groupi_n_2094));
dff csa_tree_add_14_36_groupi_retime_s1_70_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1097), .q(csa_tree_add_14_36_groupi_n_2093));
dff csa_tree_add_14_36_groupi_retime_s1_71_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_690), .q(csa_tree_add_14_36_groupi_n_2092));
dff csa_tree_add_14_36_groupi_retime_s1_72_reg (.reset(reset), .ck(clk), .d(n_2514), .q(csa_tree_add_14_36_groupi_n_2091));
dff csa_tree_add_14_36_groupi_retime_s1_73_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1067), .q(csa_tree_add_14_36_groupi_n_2090));
dff csa_tree_add_14_36_groupi_retime_s1_74_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_669), .q(csa_tree_add_14_36_groupi_n_2089));
dff csa_tree_add_14_36_groupi_retime_s1_75_reg (.reset(reset), .ck(clk), .d(n_2511), .q(csa_tree_add_14_36_groupi_n_2088));
dff csa_tree_add_14_36_groupi_retime_s1_76_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_686), .q(csa_tree_add_14_36_groupi_n_2298));
dff csa_tree_add_14_36_groupi_retime_s1_77_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_668), .q(csa_tree_add_14_36_groupi_n_2087));
dff csa_tree_add_14_36_groupi_retime_s1_78_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_630), .q(csa_tree_add_14_36_groupi_n_2086));
dff csa_tree_add_14_36_groupi_retime_s1_79_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_629), .q(csa_tree_add_14_36_groupi_n_2085));
dff csa_tree_add_14_36_groupi_retime_s1_80_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_628), .q(csa_tree_add_14_36_groupi_n_2084));
dff csa_tree_add_14_36_groupi_retime_s1_81_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_627), .q(csa_tree_add_14_36_groupi_n_2083));
dff csa_tree_add_14_36_groupi_retime_s1_82_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_626), .q(csa_tree_add_14_36_groupi_n_2082));
dff csa_tree_add_14_36_groupi_retime_s1_83_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_625), .q(csa_tree_add_14_36_groupi_n_2081));
dff csa_tree_add_14_36_groupi_retime_s1_84_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_624), .q(csa_tree_add_14_36_groupi_n_2080));
dff csa_tree_add_14_36_groupi_retime_s1_85_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_623), .q(csa_tree_add_14_36_groupi_n_2079));
dff csa_tree_add_14_36_groupi_retime_s1_86_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_622), .q(csa_tree_add_14_36_groupi_n_2078));
dff csa_tree_add_14_36_groupi_retime_s1_87_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_621), .q(csa_tree_add_14_36_groupi_n_2077));
dff csa_tree_add_14_36_groupi_retime_s1_88_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_620), .q(csa_tree_add_14_36_groupi_n_2076));
dff csa_tree_add_14_36_groupi_retime_s1_89_reg (.reset(reset), .ck(clk), .d(n_2465), .q(csa_tree_add_14_36_groupi_n_2075));
dff csa_tree_add_14_36_groupi_retime_s1_90_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_667), .q(csa_tree_add_14_36_groupi_n_2074));
dff csa_tree_add_14_36_groupi_retime_s1_91_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_763), .q(csa_tree_add_14_36_groupi_n_2073));
dff csa_tree_add_14_36_groupi_retime_s1_92_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_764), .q(csa_tree_add_14_36_groupi_n_2072));
dff csa_tree_add_14_36_groupi_retime_s1_93_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_685), .q(csa_tree_add_14_36_groupi_n_2071));
dff csa_tree_add_14_36_groupi_retime_s1_94_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_765), .q(csa_tree_add_14_36_groupi_n_2070));
dff csa_tree_add_14_36_groupi_retime_s1_95_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_766), .q(csa_tree_add_14_36_groupi_n_2069));
dff csa_tree_add_14_36_groupi_retime_s1_96_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_755), .q(csa_tree_add_14_36_groupi_n_2068));
dff csa_tree_add_14_36_groupi_retime_s1_97_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1167), .q(csa_tree_add_14_36_groupi_n_2067));
dff csa_tree_add_14_36_groupi_retime_s1_98_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_113), .q(csa_tree_add_14_36_groupi_n_2066));
dff csa_tree_add_14_36_groupi_retime_s1_99_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_500), .q(csa_tree_add_14_36_groupi_n_2065));
dff csa_tree_add_14_36_groupi_retime_s1_100_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1235), .q(csa_tree_add_14_36_groupi_n_2064));
dff csa_tree_add_14_36_groupi_retime_s1_101_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_684), .q(csa_tree_add_14_36_groupi_n_2063));
dff csa_tree_add_14_36_groupi_retime_s1_102_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_683), .q(csa_tree_add_14_36_groupi_n_2062));
dff csa_tree_add_14_36_groupi_retime_s1_103_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_701), .q(csa_tree_add_14_36_groupi_n_2061));
dff csa_tree_add_14_36_groupi_retime_s1_104_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_697), .q(csa_tree_add_14_36_groupi_n_2060));
dff csa_tree_add_14_36_groupi_retime_s1_105_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_681), .q(csa_tree_add_14_36_groupi_n_2059));
dff csa_tree_add_14_36_groupi_retime_s1_106_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_680), .q(csa_tree_add_14_36_groupi_n_2058));
dff csa_tree_add_14_36_groupi_retime_s1_107_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_679), .q(csa_tree_add_14_36_groupi_n_2057));
dff csa_tree_add_14_36_groupi_retime_s1_108_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_678), .q(csa_tree_add_14_36_groupi_n_2056));
dff csa_tree_add_14_36_groupi_retime_s1_109_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_677), .q(csa_tree_add_14_36_groupi_n_2055));
dff csa_tree_add_14_36_groupi_retime_s1_110_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_676), .q(csa_tree_add_14_36_groupi_n_2054));
dff csa_tree_add_14_36_groupi_retime_s1_111_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_675), .q(csa_tree_add_14_36_groupi_n_2053));
dff csa_tree_add_14_36_groupi_retime_s1_112_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_688), .q(csa_tree_add_14_36_groupi_n_2052));
dff csa_tree_add_14_36_groupi_retime_s1_113_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_499), .q(csa_tree_add_14_36_groupi_n_2051));
dff csa_tree_add_14_36_groupi_retime_s1_114_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_767), .q(csa_tree_add_14_36_groupi_n_2050));
dff csa_tree_add_14_36_groupi_retime_s1_115_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_768), .q(csa_tree_add_14_36_groupi_n_2049));
dff csa_tree_add_14_36_groupi_retime_s1_116_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1165), .q(csa_tree_add_14_36_groupi_n_2048));
dff csa_tree_add_14_36_groupi_retime_s1_117_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_699), .q(csa_tree_add_14_36_groupi_n_2047));
dff csa_tree_add_14_36_groupi_retime_s1_118_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1119), .q(csa_tree_add_14_36_groupi_n_2046));
dff csa_tree_add_14_36_groupi_retime_s1_119_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_769), .q(csa_tree_add_14_36_groupi_n_2045));
dff csa_tree_add_14_36_groupi_retime_s1_120_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_754), .q(csa_tree_add_14_36_groupi_n_2044));
dff csa_tree_add_14_36_groupi_retime_s1_121_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_756), .q(csa_tree_add_14_36_groupi_n_2043));
dff csa_tree_add_14_36_groupi_retime_s1_122_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_682), .q(csa_tree_add_14_36_groupi_n_2042));
dff csa_tree_add_14_36_groupi_retime_s1_123_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_666), .q(csa_tree_add_14_36_groupi_n_2041));
dff csa_tree_add_14_36_groupi_retime_s1_124_reg (.reset(reset), .ck(clk), .d(n_2459), .q(csa_tree_add_14_36_groupi_n_2040));
dff csa_tree_add_14_36_groupi_retime_s1_125_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_757), .q(csa_tree_add_14_36_groupi_n_2039));
dff csa_tree_add_14_36_groupi_retime_s1_126_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_674), .q(csa_tree_add_14_36_groupi_n_2038));
dff csa_tree_add_14_36_groupi_retime_s1_127_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1163), .q(csa_tree_add_14_36_groupi_n_2037));
dff csa_tree_add_14_36_groupi_retime_s1_128_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_240), .q(csa_tree_add_14_36_groupi_n_2036));
dff csa_tree_add_14_36_groupi_retime_s1_129_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_114), .q(csa_tree_add_14_36_groupi_n_2035));
dff csa_tree_add_14_36_groupi_retime_s1_130_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_116), .q(csa_tree_add_14_36_groupi_n_2034));
dff csa_tree_add_14_36_groupi_retime_s1_131_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_93), .q(csa_tree_add_14_36_groupi_n_2033));
dff csa_tree_add_14_36_groupi_retime_s1_132_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_673), .q(csa_tree_add_14_36_groupi_n_2032));
dff csa_tree_add_14_36_groupi_retime_s1_133_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_692), .q(csa_tree_add_14_36_groupi_n_2031));
dff csa_tree_add_14_36_groupi_retime_s1_134_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_495), .q(csa_tree_add_14_36_groupi_n_2030));
dff csa_tree_add_14_36_groupi_retime_s1_135_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_633), .q(csa_tree_add_14_36_groupi_n_2029));
dff csa_tree_add_14_36_groupi_retime_s1_136_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_90), .q(csa_tree_add_14_36_groupi_n_2028));
dff csa_tree_add_14_36_groupi_retime_s1_137_reg (.reset(reset), .ck(clk), .d(n_2440), .q(csa_tree_add_14_36_groupi_n_2027));
dff csa_tree_add_14_36_groupi_retime_s1_138_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_330), .q(csa_tree_add_14_36_groupi_n_2026));
dff csa_tree_add_14_36_groupi_retime_s1_139_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_770), .q(csa_tree_add_14_36_groupi_n_2025));
dff csa_tree_add_14_36_groupi_retime_s1_140_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_771), .q(csa_tree_add_14_36_groupi_n_2024));
dff csa_tree_add_14_36_groupi_retime_s1_141_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_115), .q(csa_tree_add_14_36_groupi_n_2297));
dff csa_tree_add_14_36_groupi_retime_s1_142_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_663), .q(csa_tree_add_14_36_groupi_n_2023));
dff csa_tree_add_14_36_groupi_retime_s2_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_48), .q(csa_tree_add_14_36_groupi_n_2174));
dff csa_tree_add_14_36_groupi_retime_s2_3_reg (.reset(reset), .ck(clk), .d(n_2570), .q(csa_tree_add_14_36_groupi_n_2169));
dff csa_tree_add_14_36_groupi_retime_s2_4_reg (.reset(reset), .ck(clk), .d(n_2569), .q(csa_tree_add_14_36_groupi_n_2168));
dff csa_tree_add_14_36_groupi_retime_s2_5_reg (.reset(reset), .ck(clk), .d(n_2437), .q(csa_tree_add_14_36_groupi_n_2166));
dff csa_tree_add_14_36_groupi_retime_s2_9_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_2142), .q(csa_tree_add_14_36_groupi_n_2141));
dff csa_tree_add_14_36_groupi_retime_s2_10_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_2139), .q(csa_tree_add_14_36_groupi_n_2138));
dff csa_tree_add_14_36_groupi_retime_s2_12_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_2098), .q(csa_tree_add_14_36_groupi_n_2097));
dff csa_tree_add_14_36_groupi_retime_s3_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1914), .q(csa_tree_add_14_36_groupi_n_2259));
dff csa_tree_add_14_36_groupi_retime_s5_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1572), .q(csa_tree_add_14_36_groupi_n_2179));
dff csa_tree_add_14_36_groupi_retime_s5_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1530), .q(csa_tree_add_14_36_groupi_n_2178));
dff csa_tree_add_14_36_groupi_retime_s5_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1436), .q(csa_tree_add_14_36_groupi_n_2176));
dff csa_tree_add_14_36_groupi_retime_s5_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1556), .q(csa_tree_add_14_36_groupi_n_2175));
dff csa_tree_add_14_36_groupi_retime_s5_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1688), .q(csa_tree_add_14_36_groupi_n_2173));
dff csa_tree_add_14_36_groupi_retime_s5_7_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1615), .q(csa_tree_add_14_36_groupi_n_2172));
dff csa_tree_add_14_36_groupi_retime_s5_8_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1767), .q(csa_tree_add_14_36_groupi_n_2171));
dff csa_tree_add_14_36_groupi_retime_s5_9_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1507), .q(csa_tree_add_14_36_groupi_n_2170));
dff csa_tree_add_14_36_groupi_retime_s5_10_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1614), .q(csa_tree_add_14_36_groupi_n_2165));
dff csa_tree_add_14_36_groupi_retime_s5_11_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1613), .q(csa_tree_add_14_36_groupi_n_2163));
dff csa_tree_add_14_36_groupi_retime_s5_12_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1687), .q(csa_tree_add_14_36_groupi_n_2162));
dff csa_tree_add_14_36_groupi_retime_s5_13_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1650), .q(csa_tree_add_14_36_groupi_n_2161));
dff csa_tree_add_14_36_groupi_retime_s5_14_reg (.reset(reset), .ck(clk), .d(n_2436), .q(csa_tree_add_14_36_groupi_n_2160));
dff csa_tree_add_14_36_groupi_retime_s5_15_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1357), .q(csa_tree_add_14_36_groupi_n_2159));
dff csa_tree_add_14_36_groupi_retime_s6_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1960), .q(csa_tree_add_14_36_groupi_n_2258));
dff csa_tree_add_14_36_groupi_retime_s6_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1833), .q(csa_tree_add_14_36_groupi_n_2177));
dff csa_tree_add_14_36_groupi_retime_s8_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1677), .q(csa_tree_add_14_36_groupi_n_2186));
dff csa_tree_add_14_36_groupi_retime_s8_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1623), .q(csa_tree_add_14_36_groupi_n_2185));
dff csa_tree_add_14_36_groupi_retime_s8_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1528), .q(csa_tree_add_14_36_groupi_n_2184));
dff csa_tree_add_14_36_groupi_retime_s8_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1532), .q(csa_tree_add_14_36_groupi_n_2183));
dff csa_tree_add_14_36_groupi_retime_s8_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1585), .q(csa_tree_add_14_36_groupi_n_2182));
dff csa_tree_add_14_36_groupi_retime_s8_7_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1565), .q(csa_tree_add_14_36_groupi_n_2181));
dff csa_tree_add_14_36_groupi_retime_s8_8_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1590), .q(csa_tree_add_14_36_groupi_n_2180));
dff csa_tree_add_14_36_groupi_retime_s8_9_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1589), .q(csa_tree_add_14_36_groupi_n_2164));
dff csa_tree_add_14_36_groupi_retime_s9_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1886), .q(csa_tree_add_14_36_groupi_n_2257));
dff csa_tree_add_14_36_groupi_retime_s9_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1855), .q(csa_tree_add_14_36_groupi_n_2188));
dff csa_tree_add_14_36_groupi_retime_s9_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1961), .q(csa_tree_add_14_36_groupi_n_2187));
dff csa_tree_add_14_36_groupi_retime_s11_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1529), .q(csa_tree_add_14_36_groupi_n_2256));
dff csa_tree_add_14_36_groupi_retime_s11_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1534), .q(csa_tree_add_14_36_groupi_n_2196));
dff csa_tree_add_14_36_groupi_retime_s11_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1554), .q(csa_tree_add_14_36_groupi_n_2193));
dff csa_tree_add_14_36_groupi_retime_s11_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1667), .q(csa_tree_add_14_36_groupi_n_2192));
dff csa_tree_add_14_36_groupi_retime_s11_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1678), .q(csa_tree_add_14_36_groupi_n_2191));
dff csa_tree_add_14_36_groupi_retime_s11_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1649), .q(csa_tree_add_14_36_groupi_n_2189));
dff csa_tree_add_14_36_groupi_retime_s12_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_52), .q(csa_tree_add_14_36_groupi_n_2199));
dff csa_tree_add_14_36_groupi_retime_s12_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1904), .q(csa_tree_add_14_36_groupi_n_2198));
dff csa_tree_add_14_36_groupi_retime_s12_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1881), .q(csa_tree_add_14_36_groupi_n_2197));
dff csa_tree_add_14_36_groupi_retime_s12_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1891), .q(csa_tree_add_14_36_groupi_n_2195));
dff csa_tree_add_14_36_groupi_retime_s12_7_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1964), .q(csa_tree_add_14_36_groupi_n_2194));
dff csa_tree_add_14_36_groupi_retime_s12_8_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1873), .q(csa_tree_add_14_36_groupi_n_2190));
dff csa_tree_add_14_36_groupi_retime_s14_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1435), .q(csa_tree_add_14_36_groupi_n_2255));
dff csa_tree_add_14_36_groupi_retime_s14_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1648), .q(csa_tree_add_14_36_groupi_n_2205));
dff csa_tree_add_14_36_groupi_retime_s14_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1587), .q(csa_tree_add_14_36_groupi_n_2204));
dff csa_tree_add_14_36_groupi_retime_s14_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1714), .q(csa_tree_add_14_36_groupi_n_2203));
dff csa_tree_add_14_36_groupi_retime_s14_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1531), .q(csa_tree_add_14_36_groupi_n_2202));
dff csa_tree_add_14_36_groupi_retime_s14_7_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1557), .q(csa_tree_add_14_36_groupi_n_2201));
dff csa_tree_add_14_36_groupi_retime_s14_8_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1668), .q(csa_tree_add_14_36_groupi_n_2200));
dff csa_tree_add_14_36_groupi_retime_s15_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1876), .q(csa_tree_add_14_36_groupi_n_2206));
dff csa_tree_add_14_36_groupi_retime_s17_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1562), .q(csa_tree_add_14_36_groupi_n_2254));
dff csa_tree_add_14_36_groupi_retime_s17_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1440), .q(csa_tree_add_14_36_groupi_n_2216));
dff csa_tree_add_14_36_groupi_retime_s17_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1591), .q(csa_tree_add_14_36_groupi_n_2209));
dff csa_tree_add_14_36_groupi_retime_s17_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1486), .q(csa_tree_add_14_36_groupi_n_2208));
dff csa_tree_add_14_36_groupi_retime_s17_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1510), .q(csa_tree_add_14_36_groupi_n_2207));
dff csa_tree_add_14_36_groupi_retime_s18_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1894), .q(csa_tree_add_14_36_groupi_n_2220));
dff csa_tree_add_14_36_groupi_retime_s18_3_reg (.reset(reset), .ck(clk), .d(n_2505), .q(csa_tree_add_14_36_groupi_n_2217));
dff csa_tree_add_14_36_groupi_retime_s18_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1923), .q(csa_tree_add_14_36_groupi_n_2215));
dff csa_tree_add_14_36_groupi_retime_s18_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1925), .q(csa_tree_add_14_36_groupi_n_2212));
dff csa_tree_add_14_36_groupi_retime_s18_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1892), .q(csa_tree_add_14_36_groupi_n_2211));
dff csa_tree_add_14_36_groupi_retime_s18_7_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1897), .q(csa_tree_add_14_36_groupi_n_2210));
dff csa_tree_add_14_36_groupi_retime_s20_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1533), .q(csa_tree_add_14_36_groupi_n_2253));
dff csa_tree_add_14_36_groupi_retime_s20_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1535), .q(csa_tree_add_14_36_groupi_n_2226));
dff csa_tree_add_14_36_groupi_retime_s20_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1679), .q(csa_tree_add_14_36_groupi_n_2225));
dff csa_tree_add_14_36_groupi_retime_s20_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1653), .q(csa_tree_add_14_36_groupi_n_2224));
dff csa_tree_add_14_36_groupi_retime_s20_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1487), .q(csa_tree_add_14_36_groupi_n_2223));
dff csa_tree_add_14_36_groupi_retime_s20_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1685), .q(csa_tree_add_14_36_groupi_n_2222));
dff csa_tree_add_14_36_groupi_retime_s20_8_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1683), .q(csa_tree_add_14_36_groupi_n_2219));
dff csa_tree_add_14_36_groupi_retime_s20_9_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1684), .q(csa_tree_add_14_36_groupi_n_2218));
dff csa_tree_add_14_36_groupi_retime_s20_10_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1802), .q(csa_tree_add_14_36_groupi_n_2214));
dff csa_tree_add_14_36_groupi_retime_s20_11_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1742), .q(csa_tree_add_14_36_groupi_n_2213));
dff csa_tree_add_14_36_groupi_retime_s21_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1866), .q(csa_tree_add_14_36_groupi_n_2228));
dff csa_tree_add_14_36_groupi_retime_s21_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_53), .q(csa_tree_add_14_36_groupi_n_2227));
dff csa_tree_add_14_36_groupi_retime_s21_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1890), .q(csa_tree_add_14_36_groupi_n_2221));
dff csa_tree_add_14_36_groupi_retime_s23_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1652), .q(csa_tree_add_14_36_groupi_n_2229));
dff csa_tree_add_14_36_groupi_retime_s24_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1863), .q(csa_tree_add_14_36_groupi_n_2252));
dff csa_tree_add_14_36_groupi_retime_s24_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1868), .q(csa_tree_add_14_36_groupi_n_2251));
dff csa_tree_add_14_36_groupi_retime_s24_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1848), .q(csa_tree_add_14_36_groupi_n_2231));
dff csa_tree_add_14_36_groupi_retime_s24_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1899), .q(csa_tree_add_14_36_groupi_n_2230));
dff csa_tree_add_14_36_groupi_retime_s26_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1686), .q(csa_tree_add_14_36_groupi_n_2249));
dff csa_tree_add_14_36_groupi_retime_s26_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1607), .q(csa_tree_add_14_36_groupi_n_2246));
dff csa_tree_add_14_36_groupi_retime_s26_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1657), .q(csa_tree_add_14_36_groupi_n_2244));
dff csa_tree_add_14_36_groupi_retime_s26_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1584), .q(csa_tree_add_14_36_groupi_n_2241));
dff csa_tree_add_14_36_groupi_retime_s26_8_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1563), .q(csa_tree_add_14_36_groupi_n_2238));
dff csa_tree_add_14_36_groupi_retime_s26_9_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1619), .q(csa_tree_add_14_36_groupi_n_2237));
dff csa_tree_add_14_36_groupi_retime_s26_10_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1715), .q(csa_tree_add_14_36_groupi_n_2236));
dff csa_tree_add_14_36_groupi_retime_s26_11_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1656), .q(csa_tree_add_14_36_groupi_n_2232));
dff csa_tree_add_14_36_groupi_retime_s27_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_2313), .q(csa_tree_add_14_36_groupi_n_2250));
dff csa_tree_add_14_36_groupi_retime_s27_2_reg (.reset(reset), .ck(clk), .d(n_2485), .q(csa_tree_add_14_36_groupi_n_2248));
dff csa_tree_add_14_36_groupi_retime_s27_3_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1744), .q(csa_tree_add_14_36_groupi_n_2247));
dff csa_tree_add_14_36_groupi_retime_s27_4_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_2246), .q(csa_tree_add_14_36_groupi_n_2245));
dff csa_tree_add_14_36_groupi_retime_s27_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1717), .q(csa_tree_add_14_36_groupi_n_2243));
dff csa_tree_add_14_36_groupi_retime_s27_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1733), .q(csa_tree_add_14_36_groupi_n_2242));
dff csa_tree_add_14_36_groupi_retime_s27_7_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_2312), .q(csa_tree_add_14_36_groupi_n_2240));
dff csa_tree_add_14_36_groupi_retime_s27_9_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1743), .q(csa_tree_add_14_36_groupi_n_2239));
dff csa_tree_add_14_36_groupi_retime_s27_10_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1792), .q(csa_tree_add_14_36_groupi_n_2235));
dff csa_tree_add_14_36_groupi_retime_s27_11_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1929), .q(csa_tree_add_14_36_groupi_n_2234));
dff csa_tree_add_14_36_groupi_retime_s27_12_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_1815), .q(csa_tree_add_14_36_groupi_n_2233));
xor2 csa_tree_add_14_36_groupi_g50786__8780 (.a(csa_tree_add_14_36_groupi_n_2020), .b(csa_tree_add_14_36_groupi_n_1812), .y(result_0__28_));
xor2 csa_tree_add_14_36_groupi_g50787__4296 (.a(csa_tree_add_14_36_groupi_n_2014), .b(csa_tree_add_14_36_groupi_n_2231), .y(result_0__25_));
xor2 csa_tree_add_14_36_groupi_g50788__3772 (.a(csa_tree_add_14_36_groupi_n_2019), .b(csa_tree_add_14_36_groupi_n_1730), .y(result_0__30_));
xor2 csa_tree_add_14_36_groupi_g50789__1474 (.a(csa_tree_add_14_36_groupi_n_2018), .b(csa_tree_add_14_36_groupi_n_1827), .y(result_0__27_));
xor2 csa_tree_add_14_36_groupi_g50790__4547 (.a(csa_tree_add_14_36_groupi_n_2017), .b(csa_tree_add_14_36_groupi_n_2233), .y(result_0__26_));
nand2 csa_tree_add_14_36_groupi_g50791__9682 (.a(csa_tree_add_14_36_groupi_n_2022), .b(csa_tree_add_14_36_groupi_n_1996), .y(result_0__29_));
nand2 csa_tree_add_14_36_groupi_g50792__2683 (.a(csa_tree_add_14_36_groupi_n_2016), .b(csa_tree_add_14_36_groupi_n_2015), .y(result_0__31_));
inv csa_tree_add_14_36_groupi_g50793 (.a(csa_tree_add_14_36_groupi_n_2021), .y(csa_tree_add_14_36_groupi_n_2022));
nand2 csa_tree_add_14_36_groupi_g50794__1309 (.a(csa_tree_add_14_36_groupi_n_2007), .b(csa_tree_add_14_36_groupi_n_2009), .y(csa_tree_add_14_36_groupi_n_2021));
nor2 csa_tree_add_14_36_groupi_g50795__6877 (.a(csa_tree_add_14_36_groupi_n_2006), .b(csa_tree_add_14_36_groupi_n_1965), .y(csa_tree_add_14_36_groupi_n_2020));
nand2 csa_tree_add_14_36_groupi_g50796__2900 (.a(csa_tree_add_14_36_groupi_n_2013), .b(csa_tree_add_14_36_groupi_n_1974), .y(csa_tree_add_14_36_groupi_n_2019));
nor2 csa_tree_add_14_36_groupi_g50797__2391 (.a(csa_tree_add_14_36_groupi_n_2011), .b(csa_tree_add_14_36_groupi_n_2234), .y(csa_tree_add_14_36_groupi_n_2018));
nand2 csa_tree_add_14_36_groupi_g50798__7675 (.a(csa_tree_add_14_36_groupi_n_2008), .b(csa_tree_add_14_36_groupi_n_2230), .y(csa_tree_add_14_36_groupi_n_2017));
nand2 csa_tree_add_14_36_groupi_g50799__7118 (.a(csa_tree_add_14_36_groupi_n_2013), .b(csa_tree_add_14_36_groupi_n_1985), .y(csa_tree_add_14_36_groupi_n_2016));
nor2 csa_tree_add_14_36_groupi_g50800__8757 (.a(csa_tree_add_14_36_groupi_n_2010), .b(csa_tree_add_14_36_groupi_n_1990), .y(csa_tree_add_14_36_groupi_n_2015));
xor2 csa_tree_add_14_36_groupi_g50801__1786 (.a(csa_tree_add_14_36_groupi_n_2003), .b(csa_tree_add_14_36_groupi_n_1934), .y(result_0__21_));
xor2 csa_tree_add_14_36_groupi_g50802__5953 (.a(csa_tree_add_14_36_groupi_n_2005), .b(csa_tree_add_14_36_groupi_n_1889), .y(result_0__24_));
xor2 csa_tree_add_14_36_groupi_g50803__5703 (.a(csa_tree_add_14_36_groupi_n_2002), .b(csa_tree_add_14_36_groupi_n_1910), .y(result_0__23_));
nor2 csa_tree_add_14_36_groupi_g50804__7114 (.a(csa_tree_add_14_36_groupi_n_2012), .b(csa_tree_add_14_36_groupi_n_84), .y(csa_tree_add_14_36_groupi_n_2014));
nor2 csa_tree_add_14_36_groupi_g50805__5266 (.a(csa_tree_add_14_36_groupi_n_2005), .b(csa_tree_add_14_36_groupi_n_2252), .y(csa_tree_add_14_36_groupi_n_2012));
nor2 csa_tree_add_14_36_groupi_g50806__2250 (.a(csa_tree_add_14_36_groupi_n_2005), .b(csa_tree_add_14_36_groupi_n_1917), .y(csa_tree_add_14_36_groupi_n_2011));
nor2 csa_tree_add_14_36_groupi_g50807__6083 (.a(csa_tree_add_14_36_groupi_n_2005), .b(csa_tree_add_14_36_groupi_n_1956), .y(csa_tree_add_14_36_groupi_n_2010));
nand2 csa_tree_add_14_36_groupi_g50808__2703 (.a(csa_tree_add_14_36_groupi_n_2004), .b(csa_tree_add_14_36_groupi_n_1945), .y(csa_tree_add_14_36_groupi_n_2013));
nand2 csa_tree_add_14_36_groupi_g50809__5795 (.a(csa_tree_add_14_36_groupi_n_2005), .b(csa_tree_add_14_36_groupi_n_1978), .y(csa_tree_add_14_36_groupi_n_2009));
nand2 csa_tree_add_14_36_groupi_g50810__7344 (.a(csa_tree_add_14_36_groupi_n_2004), .b(csa_tree_add_14_36_groupi_n_2251), .y(csa_tree_add_14_36_groupi_n_2008));
nand2 csa_tree_add_14_36_groupi_g50811__1840 (.a(csa_tree_add_14_36_groupi_n_2004), .b(csa_tree_add_14_36_groupi_n_1947), .y(csa_tree_add_14_36_groupi_n_2007));
nor2 csa_tree_add_14_36_groupi_g50812__5019 (.a(csa_tree_add_14_36_groupi_n_2005), .b(csa_tree_add_14_36_groupi_n_1932), .y(csa_tree_add_14_36_groupi_n_2006));
inv csa_tree_add_14_36_groupi_g50813 (.a(csa_tree_add_14_36_groupi_n_2005), .y(csa_tree_add_14_36_groupi_n_2004));
nand2 csa_tree_add_14_36_groupi_g50814__1857 (.a(csa_tree_add_14_36_groupi_n_2001), .b(csa_tree_add_14_36_groupi_n_2215), .y(csa_tree_add_14_36_groupi_n_2003));
nand2 csa_tree_add_14_36_groupi_g50815__9906 (.a(csa_tree_add_14_36_groupi_n_2000), .b(csa_tree_add_14_36_groupi_n_2221), .y(csa_tree_add_14_36_groupi_n_2002));
nor2 csa_tree_add_14_36_groupi_g50816__8780 (.a(csa_tree_add_14_36_groupi_n_1998), .b(csa_tree_add_14_36_groupi_n_1967), .y(csa_tree_add_14_36_groupi_n_2005));
xor2 csa_tree_add_14_36_groupi_g50817__4296 (.a(csa_tree_add_14_36_groupi_n_1994), .b(csa_tree_add_14_36_groupi_n_1946), .y(result_0__20_));
xor2 csa_tree_add_14_36_groupi_g50818__3772 (.a(csa_tree_add_14_36_groupi_n_1997), .b(csa_tree_add_14_36_groupi_n_1927), .y(result_0__22_));
xor2 csa_tree_add_14_36_groupi_g50819__1474 (.a(csa_tree_add_14_36_groupi_n_1995), .b(csa_tree_add_14_36_groupi_n_1926), .y(result_0__19_));
nand2 csa_tree_add_14_36_groupi_g50820__4547 (.a(csa_tree_add_14_36_groupi_n_1993), .b(csa_tree_add_14_36_groupi_n_2212), .y(csa_tree_add_14_36_groupi_n_2001));
inv csa_tree_add_14_36_groupi_g50821 (.a(csa_tree_add_14_36_groupi_n_1999), .y(csa_tree_add_14_36_groupi_n_2000));
nor2 csa_tree_add_14_36_groupi_g50822__9682 (.a(csa_tree_add_14_36_groupi_n_1997), .b(csa_tree_add_14_36_groupi_n_2316), .y(csa_tree_add_14_36_groupi_n_1999));
nor2 csa_tree_add_14_36_groupi_g50823__2683 (.a(csa_tree_add_14_36_groupi_n_1994), .b(csa_tree_add_14_36_groupi_n_1952), .y(csa_tree_add_14_36_groupi_n_1998));
nor2 csa_tree_add_14_36_groupi_g50824__1309 (.a(csa_tree_add_14_36_groupi_n_1991), .b(csa_tree_add_14_36_groupi_n_1980), .y(csa_tree_add_14_36_groupi_n_1996));
nand2 csa_tree_add_14_36_groupi_g50825__6877 (.a(csa_tree_add_14_36_groupi_n_1992), .b(csa_tree_add_14_36_groupi_n_2317), .y(csa_tree_add_14_36_groupi_n_1995));
nor2 csa_tree_add_14_36_groupi_g50826__2900 (.a(csa_tree_add_14_36_groupi_n_1963), .b(csa_tree_add_14_36_groupi_n_1989), .y(csa_tree_add_14_36_groupi_n_1997));
inv csa_tree_add_14_36_groupi_g50827 (.a(csa_tree_add_14_36_groupi_n_1993), .y(csa_tree_add_14_36_groupi_n_1994));
xor2 csa_tree_add_14_36_groupi_g50828__2391 (.a(csa_tree_add_14_36_groupi_n_1982), .b(csa_tree_add_14_36_groupi_n_2305), .y(result_0__17_));
xor2 csa_tree_add_14_36_groupi_g50829__7675 (.a(csa_tree_add_14_36_groupi_n_1986), .b(csa_tree_add_14_36_groupi_n_1921), .y(result_0__18_));
xor2 csa_tree_add_14_36_groupi_g50830__7118 (.a(csa_tree_add_14_36_groupi_n_1981), .b(csa_tree_add_14_36_groupi_n_2195), .y(result_0__15_));
nand2 csa_tree_add_14_36_groupi_g50831__8757 (.a(csa_tree_add_14_36_groupi_n_1988), .b(csa_tree_add_14_36_groupi_n_1944), .y(csa_tree_add_14_36_groupi_n_1993));
nand2 csa_tree_add_14_36_groupi_g50832__1786 (.a(csa_tree_add_14_36_groupi_n_1987), .b(csa_tree_add_14_36_groupi_n_2206), .y(csa_tree_add_14_36_groupi_n_1992));
nand2 csa_tree_add_14_36_groupi_g50833__5953 (.a(csa_tree_add_14_36_groupi_n_1983), .b(csa_tree_add_14_36_groupi_n_1979), .y(csa_tree_add_14_36_groupi_n_1991));
nand2 csa_tree_add_14_36_groupi_g50834__5703 (.a(csa_tree_add_14_36_groupi_n_1984), .b(csa_tree_add_14_36_groupi_n_1790), .y(csa_tree_add_14_36_groupi_n_1990));
nor2 csa_tree_add_14_36_groupi_g50835__7114 (.a(csa_tree_add_14_36_groupi_n_1953), .b(csa_tree_add_14_36_groupi_n_1986), .y(csa_tree_add_14_36_groupi_n_1989));
nand2 csa_tree_add_14_36_groupi_g50836__5266 (.a(csa_tree_add_14_36_groupi_n_1987), .b(csa_tree_add_14_36_groupi_n_1933), .y(csa_tree_add_14_36_groupi_n_1988));
inv csa_tree_add_14_36_groupi_g50837 (.a(csa_tree_add_14_36_groupi_n_1987), .y(csa_tree_add_14_36_groupi_n_1986));
nor2 csa_tree_add_14_36_groupi_g50838__2250 (.a(csa_tree_add_14_36_groupi_n_1975), .b(csa_tree_add_14_36_groupi_n_1735), .y(csa_tree_add_14_36_groupi_n_1985));
nand2 csa_tree_add_14_36_groupi_g50839__6083 (.a(csa_tree_add_14_36_groupi_n_1975), .b(csa_tree_add_14_36_groupi_n_313), .y(csa_tree_add_14_36_groupi_n_1984));
nand2 csa_tree_add_14_36_groupi_g50840__2703 (.a(csa_tree_add_14_36_groupi_n_1972), .b(csa_tree_add_14_36_groupi_n_1814), .y(csa_tree_add_14_36_groupi_n_1983));
nand2 csa_tree_add_14_36_groupi_g50841__5795 (.a(csa_tree_add_14_36_groupi_n_1977), .b(csa_tree_add_14_36_groupi_n_2318), .y(csa_tree_add_14_36_groupi_n_1982));
nor2 csa_tree_add_14_36_groupi_g50842__7344 (.a(csa_tree_add_14_36_groupi_n_1971), .b(csa_tree_add_14_36_groupi_n_2257), .y(csa_tree_add_14_36_groupi_n_1981));
nand2 csa_tree_add_14_36_groupi_g50843__1840 (.a(csa_tree_add_14_36_groupi_n_1976), .b(csa_tree_add_14_36_groupi_n_2198), .y(csa_tree_add_14_36_groupi_n_1987));
nor2 csa_tree_add_14_36_groupi_g50844__5019 (.a(csa_tree_add_14_36_groupi_n_1972), .b(csa_tree_add_14_36_groupi_n_1805), .y(csa_tree_add_14_36_groupi_n_1980));
nand2 csa_tree_add_14_36_groupi_g50845__1857 (.a(csa_tree_add_14_36_groupi_n_1972), .b(csa_tree_add_14_36_groupi_n_1939), .y(csa_tree_add_14_36_groupi_n_1979));
nor2 csa_tree_add_14_36_groupi_g50846__9906 (.a(csa_tree_add_14_36_groupi_n_1973), .b(csa_tree_add_14_36_groupi_n_1806), .y(csa_tree_add_14_36_groupi_n_1978));
xor2 csa_tree_add_14_36_groupi_g50847__8780 (.a(csa_tree_add_14_36_groupi_n_1907), .b(csa_tree_add_14_36_groupi_n_2194), .y(result_0__16_));
xor2 csa_tree_add_14_36_groupi_g50848__4296 (.a(csa_tree_add_14_36_groupi_n_1909), .b(csa_tree_add_14_36_groupi_n_2187), .y(result_0__14_));
xor2 csa_tree_add_14_36_groupi_g50849__3772 (.a(csa_tree_add_14_36_groupi_n_2258), .b(csa_tree_add_14_36_groupi_n_2188), .y(result_0__13_));
nand2 csa_tree_add_14_36_groupi_g50850__1474 (.a(csa_tree_add_14_36_groupi_n_2199), .b(csa_tree_add_14_36_groupi_n_2194), .y(csa_tree_add_14_36_groupi_n_1977));
nand2 csa_tree_add_14_36_groupi_g50851__4547 (.a(csa_tree_add_14_36_groupi_n_2197), .b(csa_tree_add_14_36_groupi_n_2194), .y(csa_tree_add_14_36_groupi_n_1976));
inv csa_tree_add_14_36_groupi_g50852 (.a(csa_tree_add_14_36_groupi_n_1974), .y(csa_tree_add_14_36_groupi_n_1975));
inv csa_tree_add_14_36_groupi_g50853 (.a(csa_tree_add_14_36_groupi_n_1972), .y(csa_tree_add_14_36_groupi_n_1973));
nor2 csa_tree_add_14_36_groupi_g50854__9682 (.a(csa_tree_add_14_36_groupi_n_2187), .b(csa_tree_add_14_36_groupi_n_1908), .y(csa_tree_add_14_36_groupi_n_1971));
nor2 csa_tree_add_14_36_groupi_g50855__2683 (.a(csa_tree_add_14_36_groupi_n_1968), .b(csa_tree_add_14_36_groupi_n_1857), .y(csa_tree_add_14_36_groupi_n_1974));
nor2 csa_tree_add_14_36_groupi_g50856__1309 (.a(csa_tree_add_14_36_groupi_n_1970), .b(csa_tree_add_14_36_groupi_n_2248), .y(csa_tree_add_14_36_groupi_n_1972));
inv csa_tree_add_14_36_groupi_g50860 (.a(csa_tree_add_14_36_groupi_n_1969), .y(csa_tree_add_14_36_groupi_n_1970));
nand2 csa_tree_add_14_36_groupi_g50861__6877 (.a(csa_tree_add_14_36_groupi_n_1965), .b(csa_tree_add_14_36_groupi_n_2247), .y(csa_tree_add_14_36_groupi_n_1969));
nor2 csa_tree_add_14_36_groupi_g50862__2900 (.a(csa_tree_add_14_36_groupi_n_1966), .b(csa_tree_add_14_36_groupi_n_1838), .y(csa_tree_add_14_36_groupi_n_1968));
nand2 csa_tree_add_14_36_groupi_g50863__2391 (.a(csa_tree_add_14_36_groupi_n_1962), .b(csa_tree_add_14_36_groupi_n_1948), .y(csa_tree_add_14_36_groupi_n_1967));
inv csa_tree_add_14_36_groupi_g50864 (.a(csa_tree_add_14_36_groupi_n_1965), .y(csa_tree_add_14_36_groupi_n_1966));
nand2 csa_tree_add_14_36_groupi_g50865__7675 (.a(csa_tree_add_14_36_groupi_n_1928), .b(csa_tree_add_14_36_groupi_n_1951), .y(csa_tree_add_14_36_groupi_n_1964));
nand2 csa_tree_add_14_36_groupi_g50866__7118 (.a(csa_tree_add_14_36_groupi_n_1950), .b(csa_tree_add_14_36_groupi_n_1958), .y(csa_tree_add_14_36_groupi_n_1963));
nand2 csa_tree_add_14_36_groupi_g50867__8757 (.a(csa_tree_add_14_36_groupi_n_1954), .b(csa_tree_add_14_36_groupi_n_2239), .y(csa_tree_add_14_36_groupi_n_1965));
nand2 csa_tree_add_14_36_groupi_g50868__1786 (.a(csa_tree_add_14_36_groupi_n_1959), .b(csa_tree_add_14_36_groupi_n_1919), .y(csa_tree_add_14_36_groupi_n_1962));
nor2 csa_tree_add_14_36_groupi_g50869__5953 (.a(csa_tree_add_14_36_groupi_n_1957), .b(csa_tree_add_14_36_groupi_n_1884), .y(csa_tree_add_14_36_groupi_n_1961));
nand2 csa_tree_add_14_36_groupi_g50870__5703 (.a(csa_tree_add_14_36_groupi_n_1955), .b(csa_tree_add_14_36_groupi_n_1776), .y(csa_tree_add_14_36_groupi_n_1960));
xor2 csa_tree_add_14_36_groupi_g50871__7114 (.a(csa_tree_add_14_36_groupi_n_1941), .b(csa_tree_add_14_36_groupi_n_1782), .y(result_0__12_));
inv csa_tree_add_14_36_groupi_g50872 (.a(csa_tree_add_14_36_groupi_n_1958), .y(csa_tree_add_14_36_groupi_n_1959));
nor2 csa_tree_add_14_36_groupi_g50873__5266 (.a(csa_tree_add_14_36_groupi_n_1941), .b(csa_tree_add_14_36_groupi_n_1860), .y(csa_tree_add_14_36_groupi_n_1957));
nand2 csa_tree_add_14_36_groupi_g50874__2250 (.a(csa_tree_add_14_36_groupi_n_1945), .b(csa_tree_add_14_36_groupi_n_313), .y(csa_tree_add_14_36_groupi_n_1956));
nand2 csa_tree_add_14_36_groupi_g50875__6083 (.a(csa_tree_add_14_36_groupi_n_1940), .b(csa_tree_add_14_36_groupi_n_1772), .y(csa_tree_add_14_36_groupi_n_1955));
nand2 csa_tree_add_14_36_groupi_g50876__2703 (.a(csa_tree_add_14_36_groupi_n_2310), .b(csa_tree_add_14_36_groupi_n_2234), .y(csa_tree_add_14_36_groupi_n_1954));
nor2 csa_tree_add_14_36_groupi_g50877__5795 (.a(csa_tree_add_14_36_groupi_n_1949), .b(csa_tree_add_14_36_groupi_n_2220), .y(csa_tree_add_14_36_groupi_n_1958));
nand2 csa_tree_add_14_36_groupi_g50878__7344 (.a(csa_tree_add_14_36_groupi_n_1933), .b(csa_tree_add_14_36_groupi_n_1942), .y(csa_tree_add_14_36_groupi_n_1953));
nand2 csa_tree_add_14_36_groupi_g50879__1840 (.a(csa_tree_add_14_36_groupi_n_1919), .b(csa_tree_add_14_36_groupi_n_1942), .y(csa_tree_add_14_36_groupi_n_1952));
nand2 csa_tree_add_14_36_groupi_g50880__5019 (.a(csa_tree_add_14_36_groupi_n_1940), .b(csa_tree_add_14_36_groupi_n_1913), .y(csa_tree_add_14_36_groupi_n_1951));
nand2 csa_tree_add_14_36_groupi_g50881__1857 (.a(csa_tree_add_14_36_groupi_n_1943), .b(csa_tree_add_14_36_groupi_n_1942), .y(csa_tree_add_14_36_groupi_n_1950));
xor2 csa_tree_add_14_36_groupi_g50882__9906 (.a(csa_tree_add_14_36_groupi_n_2177), .b(csa_tree_add_14_36_groupi_n_2259), .y(result_0__11_));
nor2 csa_tree_add_14_36_groupi_g50883__8780 (.a(csa_tree_add_14_36_groupi_n_2217), .b(csa_tree_add_14_36_groupi_n_2215), .y(csa_tree_add_14_36_groupi_n_1949));
nor2 csa_tree_add_14_36_groupi_g50884__4296 (.a(csa_tree_add_14_36_groupi_n_1936), .b(csa_tree_add_14_36_groupi_n_2228), .y(csa_tree_add_14_36_groupi_n_1948));
nor2 csa_tree_add_14_36_groupi_g50885__3772 (.a(csa_tree_add_14_36_groupi_n_1932), .b(csa_tree_add_14_36_groupi_n_1816), .y(csa_tree_add_14_36_groupi_n_1947));
nand2 csa_tree_add_14_36_groupi_g50886__1474 (.a(csa_tree_add_14_36_groupi_n_2215), .b(csa_tree_add_14_36_groupi_n_2212), .y(csa_tree_add_14_36_groupi_n_1946));
inv csa_tree_add_14_36_groupi_g50888 (.a(csa_tree_add_14_36_groupi_n_1943), .y(csa_tree_add_14_36_groupi_n_1944));
inv csa_tree_add_14_36_groupi_g50889 (.a(csa_tree_add_14_36_groupi_n_1941), .y(csa_tree_add_14_36_groupi_n_1940));
nor2 csa_tree_add_14_36_groupi_g50890__4547 (.a(csa_tree_add_14_36_groupi_n_1931), .b(csa_tree_add_14_36_groupi_n_1806), .y(csa_tree_add_14_36_groupi_n_1939));
nor2 csa_tree_add_14_36_groupi_g50891__9682 (.a(csa_tree_add_14_36_groupi_n_1932), .b(csa_tree_add_14_36_groupi_n_1838), .y(csa_tree_add_14_36_groupi_n_1945));
nand2 csa_tree_add_14_36_groupi_g50892__2683 (.a(csa_tree_add_14_36_groupi_n_1938), .b(csa_tree_add_14_36_groupi_n_2210), .y(csa_tree_add_14_36_groupi_n_1943));
nor2 csa_tree_add_14_36_groupi_g50893__1309 (.a(csa_tree_add_14_36_groupi_n_2217), .b(csa_tree_add_14_36_groupi_n_1937), .y(csa_tree_add_14_36_groupi_n_1942));
nor2 csa_tree_add_14_36_groupi_g50894__6877 (.a(csa_tree_add_14_36_groupi_n_1930), .b(csa_tree_add_14_36_groupi_n_1902), .y(csa_tree_add_14_36_groupi_n_1941));
inv csa_tree_add_14_36_groupi_g50895 (.a(csa_tree_add_14_36_groupi_n_1935), .y(csa_tree_add_14_36_groupi_n_1938));
inv csa_tree_add_14_36_groupi_g50896 (.a(csa_tree_add_14_36_groupi_n_2212), .y(csa_tree_add_14_36_groupi_n_1937));
nor2 csa_tree_add_14_36_groupi_g50897__2900 (.a(csa_tree_add_14_36_groupi_n_2227), .b(csa_tree_add_14_36_groupi_n_2221), .y(csa_tree_add_14_36_groupi_n_1936));
nor2 csa_tree_add_14_36_groupi_g50898__2391 (.a(csa_tree_add_14_36_groupi_n_2317), .b(csa_tree_add_14_36_groupi_n_2211), .y(csa_tree_add_14_36_groupi_n_1935));
nor2 csa_tree_add_14_36_groupi_g50900__7675 (.a(csa_tree_add_14_36_groupi_n_2217), .b(csa_tree_add_14_36_groupi_n_2220), .y(csa_tree_add_14_36_groupi_n_1934));
inv csa_tree_add_14_36_groupi_g50903 (.a(csa_tree_add_14_36_groupi_n_1932), .y(csa_tree_add_14_36_groupi_n_1931));
nand2 csa_tree_add_14_36_groupi_g50904__7118 (.a(csa_tree_add_14_36_groupi_n_1911), .b(csa_tree_add_14_36_groupi_n_1799), .y(csa_tree_add_14_36_groupi_n_1930));
nand2 csa_tree_add_14_36_groupi_g50905__8757 (.a(csa_tree_add_14_36_groupi_n_1920), .b(csa_tree_add_14_36_groupi_n_1796), .y(csa_tree_add_14_36_groupi_n_1929));
nor2 csa_tree_add_14_36_groupi_g50906__1786 (.a(csa_tree_add_14_36_groupi_n_1915), .b(csa_tree_add_14_36_groupi_n_1916), .y(csa_tree_add_14_36_groupi_n_1928));
nand2 csa_tree_add_14_36_groupi_g50907__5953 (.a(csa_tree_add_14_36_groupi_n_64), .b(csa_tree_add_14_36_groupi_n_2221), .y(csa_tree_add_14_36_groupi_n_1927));
nor2 csa_tree_add_14_36_groupi_g50908__5703 (.a(csa_tree_add_14_36_groupi_n_2211), .b(csa_tree_add_14_36_groupi_n_1905), .y(csa_tree_add_14_36_groupi_n_1933));
nor2 csa_tree_add_14_36_groupi_g50909__7114 (.a(csa_tree_add_14_36_groupi_n_1924), .b(csa_tree_add_14_36_groupi_n_2211), .y(csa_tree_add_14_36_groupi_n_1926));
nand2 csa_tree_add_14_36_groupi_g50910__5266 (.a(csa_tree_add_14_36_groupi_n_1918), .b(csa_tree_add_14_36_groupi_n_2310), .y(csa_tree_add_14_36_groupi_n_1932));
inv csa_tree_add_14_36_groupi_g50911 (.a(csa_tree_add_14_36_groupi_n_1922), .y(csa_tree_add_14_36_groupi_n_1925));
inv csa_tree_add_14_36_groupi_g50912 (.a(csa_tree_add_14_36_groupi_n_2210), .y(csa_tree_add_14_36_groupi_n_1924));
nand2 csa_tree_add_14_36_groupi_g50914__2250 (.a(csa_tree_add_14_36_groupi_n_1859), .b(csa_tree_add_14_36_groupi_n_1900), .y(csa_tree_add_14_36_groupi_n_1923));
nor2 csa_tree_add_14_36_groupi_g50915__6083 (.a(csa_tree_add_14_36_groupi_n_1859), .b(csa_tree_add_14_36_groupi_n_1900), .y(csa_tree_add_14_36_groupi_n_1922));
nand2 csa_tree_add_14_36_groupi_g50917__2703 (.a(csa_tree_add_14_36_groupi_n_2317), .b(csa_tree_add_14_36_groupi_n_2206), .y(csa_tree_add_14_36_groupi_n_1921));
inv csa_tree_add_14_36_groupi_g50924 (.a(csa_tree_add_14_36_groupi_n_1912), .y(csa_tree_add_14_36_groupi_n_1920));
inv csa_tree_add_14_36_groupi_g50925 (.a(csa_tree_add_14_36_groupi_n_1917), .y(csa_tree_add_14_36_groupi_n_1918));
nand2 csa_tree_add_14_36_groupi_g50926__5795 (.a(csa_tree_add_14_36_groupi_n_1895), .b(csa_tree_add_14_36_groupi_n_1888), .y(csa_tree_add_14_36_groupi_n_1916));
xor2 csa_tree_add_14_36_groupi_g50927__7344 (.a(csa_tree_add_14_36_groupi_n_1878), .b(csa_tree_add_14_36_groupi_n_1829), .y(result_0__9_));
xor2 csa_tree_add_14_36_groupi_g50928__1840 (.a(csa_tree_add_14_36_groupi_n_1883), .b(csa_tree_add_14_36_groupi_n_1786), .y(result_0__10_));
nor2 csa_tree_add_14_36_groupi_g50929__5019 (.a(csa_tree_add_14_36_groupi_n_1885), .b(csa_tree_add_14_36_groupi_n_1898), .y(csa_tree_add_14_36_groupi_n_1915));
nand2 csa_tree_add_14_36_groupi_g50930__1857 (.a(csa_tree_add_14_36_groupi_n_1903), .b(csa_tree_add_14_36_groupi_n_1773), .y(csa_tree_add_14_36_groupi_n_1914));
nor2 csa_tree_add_14_36_groupi_g50931__9906 (.a(csa_tree_add_14_36_groupi_n_1898), .b(csa_tree_add_14_36_groupi_n_1860), .y(csa_tree_add_14_36_groupi_n_1913));
nor2 csa_tree_add_14_36_groupi_g50932__8780 (.a(csa_tree_add_14_36_groupi_n_1899), .b(csa_tree_add_14_36_groupi_n_1791), .y(csa_tree_add_14_36_groupi_n_1912));
nand2 csa_tree_add_14_36_groupi_g50933__4296 (.a(csa_tree_add_14_36_groupi_n_1896), .b(csa_tree_add_14_36_groupi_n_1793), .y(csa_tree_add_14_36_groupi_n_1911));
nor2 csa_tree_add_14_36_groupi_g50934__3772 (.a(csa_tree_add_14_36_groupi_n_2316), .b(csa_tree_add_14_36_groupi_n_2227), .y(csa_tree_add_14_36_groupi_n_1919));
nor2 csa_tree_add_14_36_groupi_g50935__1474 (.a(csa_tree_add_14_36_groupi_n_2227), .b(csa_tree_add_14_36_groupi_n_2228), .y(csa_tree_add_14_36_groupi_n_1910));
nand2 csa_tree_add_14_36_groupi_g50936__4547 (.a(csa_tree_add_14_36_groupi_n_2190), .b(csa_tree_add_14_36_groupi_n_1906), .y(csa_tree_add_14_36_groupi_n_1909));
nand2 csa_tree_add_14_36_groupi_g50937__9682 (.a(csa_tree_add_14_36_groupi_n_2235), .b(csa_tree_add_14_36_groupi_n_2251), .y(csa_tree_add_14_36_groupi_n_1917));
inv csa_tree_add_14_36_groupi_g50938 (.a(csa_tree_add_14_36_groupi_n_2190), .y(csa_tree_add_14_36_groupi_n_1908));
inv csa_tree_add_14_36_groupi_g50939 (.a(csa_tree_add_14_36_groupi_n_1901), .y(csa_tree_add_14_36_groupi_n_1907));
inv csa_tree_add_14_36_groupi_g50940 (.a(csa_tree_add_14_36_groupi_n_2257), .y(csa_tree_add_14_36_groupi_n_1906));
inv csa_tree_add_14_36_groupi_g50941 (.a(csa_tree_add_14_36_groupi_n_2206), .y(csa_tree_add_14_36_groupi_n_1905));
nor2 csa_tree_add_14_36_groupi_g50942__2683 (.a(csa_tree_add_14_36_groupi_n_1879), .b(csa_tree_add_14_36_groupi_n_1850), .y(csa_tree_add_14_36_groupi_n_1904));
nand2 csa_tree_add_14_36_groupi_g50944__1309 (.a(csa_tree_add_14_36_groupi_n_1883), .b(csa_tree_add_14_36_groupi_n_1770), .y(csa_tree_add_14_36_groupi_n_1903));
nor2 csa_tree_add_14_36_groupi_g50945__6877 (.a(csa_tree_add_14_36_groupi_n_1869), .b(csa_tree_add_14_36_groupi_n_1818), .y(csa_tree_add_14_36_groupi_n_1902));
nand2 csa_tree_add_14_36_groupi_g50948__2900 (.a(csa_tree_add_14_36_groupi_n_2318), .b(csa_tree_add_14_36_groupi_n_2199), .y(csa_tree_add_14_36_groupi_n_1901));
nand2 csa_tree_add_14_36_groupi_g50953__2391 (.a(csa_tree_add_14_36_groupi_n_1826), .b(csa_tree_add_14_36_groupi_n_1870), .y(csa_tree_add_14_36_groupi_n_1897));
nand2 csa_tree_add_14_36_groupi_g50954__7675 (.a(csa_tree_add_14_36_groupi_n_1880), .b(csa_tree_add_14_36_groupi_n_1773), .y(csa_tree_add_14_36_groupi_n_1896));
nand2 csa_tree_add_14_36_groupi_g50955__7118 (.a(csa_tree_add_14_36_groupi_n_1882), .b(csa_tree_add_14_36_groupi_n_1886), .y(csa_tree_add_14_36_groupi_n_1895));
nor2 csa_tree_add_14_36_groupi_g50956__8757 (.a(csa_tree_add_14_36_groupi_n_1875), .b(csa_tree_add_14_36_groupi_n_1871), .y(csa_tree_add_14_36_groupi_n_1894));
nor2 csa_tree_add_14_36_groupi_g50958__5953 (.a(csa_tree_add_14_36_groupi_n_1826), .b(csa_tree_add_14_36_groupi_n_1870), .y(csa_tree_add_14_36_groupi_n_1892));
nand2 csa_tree_add_14_36_groupi_g50959__5703 (.a(csa_tree_add_14_36_groupi_n_1882), .b(csa_tree_add_14_36_groupi_n_1888), .y(csa_tree_add_14_36_groupi_n_1891));
nand2 csa_tree_add_14_36_groupi_g50960__7114 (.a(csa_tree_add_14_36_groupi_n_2295), .b(n_2480), .y(csa_tree_add_14_36_groupi_n_1890));
xor2 csa_tree_add_14_36_groupi_g50961__5266 (.a(csa_tree_add_14_36_groupi_n_1777), .b(csa_tree_add_14_36_groupi_n_1844), .y(csa_tree_add_14_36_groupi_n_1900));
nand2 csa_tree_add_14_36_groupi_g50962__2250 (.a(csa_tree_add_14_36_groupi_n_2315), .b(csa_tree_add_14_36_groupi_n_1887), .y(csa_tree_add_14_36_groupi_n_1889));
nor2 csa_tree_add_14_36_groupi_g50963__6083 (.a(csa_tree_add_14_36_groupi_n_1867), .b(csa_tree_add_14_36_groupi_n_1821), .y(csa_tree_add_14_36_groupi_n_1899));
nand2 csa_tree_add_14_36_groupi_g50964__2703 (.a(csa_tree_add_14_36_groupi_n_1882), .b(csa_tree_add_14_36_groupi_n_1873), .y(csa_tree_add_14_36_groupi_n_1898));
inv csa_tree_add_14_36_groupi_g50965 (.a(csa_tree_add_14_36_groupi_n_2252), .y(csa_tree_add_14_36_groupi_n_1887));
inv csa_tree_add_14_36_groupi_g50966 (.a(csa_tree_add_14_36_groupi_n_1884), .y(csa_tree_add_14_36_groupi_n_1885));
inv csa_tree_add_14_36_groupi_g50967 (.a(csa_tree_add_14_36_groupi_n_1877), .y(csa_tree_add_14_36_groupi_n_1882));
nor2 csa_tree_add_14_36_groupi_g50968__5795 (.a(csa_tree_add_14_36_groupi_n_1849), .b(csa_tree_add_14_36_groupi_n_56), .y(csa_tree_add_14_36_groupi_n_1881));
nand2 csa_tree_add_14_36_groupi_g50969__7344 (.a(csa_tree_add_14_36_groupi_n_1862), .b(csa_tree_add_14_36_groupi_n_1770), .y(csa_tree_add_14_36_groupi_n_1880));
nor2 csa_tree_add_14_36_groupi_g50970__1840 (.a(csa_tree_add_14_36_groupi_n_1849), .b(csa_tree_add_14_36_groupi_n_2410), .y(csa_tree_add_14_36_groupi_n_1879));
nand2 csa_tree_add_14_36_groupi_g50972__5019 (.a(csa_tree_add_14_36_groupi_n_1837), .b(csa_tree_add_14_36_groupi_n_1851), .y(csa_tree_add_14_36_groupi_n_1888));
nand2 csa_tree_add_14_36_groupi_g50976__1857 (.a(csa_tree_add_14_36_groupi_n_1864), .b(csa_tree_add_14_36_groupi_n_2168), .y(csa_tree_add_14_36_groupi_n_1878));
nor2 csa_tree_add_14_36_groupi_g50977__9906 (.a(csa_tree_add_14_36_groupi_n_1853), .b(csa_tree_add_14_36_groupi_n_1738), .y(csa_tree_add_14_36_groupi_n_1886));
nand2 csa_tree_add_14_36_groupi_g50978__8780 (.a(csa_tree_add_14_36_groupi_n_1858), .b(csa_tree_add_14_36_groupi_n_1842), .y(csa_tree_add_14_36_groupi_n_1884));
nand2 csa_tree_add_14_36_groupi_g50979__4296 (.a(csa_tree_add_14_36_groupi_n_1847), .b(csa_tree_add_14_36_groupi_n_1861), .y(csa_tree_add_14_36_groupi_n_1883));
nor2 csa_tree_add_14_36_groupi_g50980__3772 (.a(csa_tree_add_14_36_groupi_n_1837), .b(csa_tree_add_14_36_groupi_n_1851), .y(csa_tree_add_14_36_groupi_n_1877));
inv csa_tree_add_14_36_groupi_g50981 (.a(csa_tree_add_14_36_groupi_n_1865), .y(csa_tree_add_14_36_groupi_n_1876));
inv csa_tree_add_14_36_groupi_g50982 (.a(n_2506), .y(csa_tree_add_14_36_groupi_n_1875));
nand2 csa_tree_add_14_36_groupi_g50984__1474 (.a(csa_tree_add_14_36_groupi_n_1793), .b(csa_tree_add_14_36_groupi_n_1845), .y(csa_tree_add_14_36_groupi_n_1869));
nor2 csa_tree_add_14_36_groupi_g50986__4547 (.a(csa_tree_add_14_36_groupi_n_1863), .b(csa_tree_add_14_36_groupi_n_1820), .y(csa_tree_add_14_36_groupi_n_1868));
nor2 csa_tree_add_14_36_groupi_g50987__9682 (.a(csa_tree_add_14_36_groupi_n_1820), .b(csa_tree_add_14_36_groupi_n_2412), .y(csa_tree_add_14_36_groupi_n_1867));
nor2 csa_tree_add_14_36_groupi_g50988__2683 (.a(csa_tree_add_14_36_groupi_n_1811), .b(n_2488), .y(csa_tree_add_14_36_groupi_n_1866));
nor2 csa_tree_add_14_36_groupi_g50989__1309 (.a(csa_tree_add_14_36_groupi_n_2294), .b(csa_tree_add_14_36_groupi_n_2293), .y(csa_tree_add_14_36_groupi_n_1865));
xor2 csa_tree_add_14_36_groupi_g50990__6877 (.a(csa_tree_add_14_36_groupi_n_1828), .b(csa_tree_add_14_36_groupi_n_1704), .y(result_0__7_));
xor2 csa_tree_add_14_36_groupi_g50991__2900 (.a(csa_tree_add_14_36_groupi_n_1818), .b(csa_tree_add_14_36_groupi_n_1693), .y(result_0__8_));
nand2 csa_tree_add_14_36_groupi_g50993__7675 (.a(csa_tree_add_14_36_groupi_n_1846), .b(n_2685), .y(csa_tree_add_14_36_groupi_n_2295));
nand2 csa_tree_add_14_36_groupi_g50994__7118 (.a(csa_tree_add_14_36_groupi_n_1853), .b(csa_tree_add_14_36_groupi_n_1738), .y(csa_tree_add_14_36_groupi_n_1873));
xor2 csa_tree_add_14_36_groupi_g50995__8757 (.a(n_2681), .b(csa_tree_add_14_36_groupi_n_2214), .y(csa_tree_add_14_36_groupi_n_1871));
xor2 csa_tree_add_14_36_groupi_g50996__1786 (.a(csa_tree_add_14_36_groupi_n_50), .b(csa_tree_add_14_36_groupi_n_1690), .y(csa_tree_add_14_36_groupi_n_1870));
inv csa_tree_add_14_36_groupi_g50997 (.a(csa_tree_add_14_36_groupi_n_1856), .y(csa_tree_add_14_36_groupi_n_1864));
inv csa_tree_add_14_36_groupi_g50998 (.a(csa_tree_add_14_36_groupi_n_1861), .y(csa_tree_add_14_36_groupi_n_1862));
nand2 csa_tree_add_14_36_groupi_g50999__5953 (.a(csa_tree_add_14_36_groupi_n_1775), .b(csa_tree_add_14_36_groupi_n_1836), .y(csa_tree_add_14_36_groupi_n_1858));
nand2 csa_tree_add_14_36_groupi_g51000__5703 (.a(csa_tree_add_14_36_groupi_n_1830), .b(csa_tree_add_14_36_groupi_n_2243), .y(csa_tree_add_14_36_groupi_n_1857));
nor2 csa_tree_add_14_36_groupi_g51001__7114 (.a(csa_tree_add_14_36_groupi_n_1818), .b(csa_tree_add_14_36_groupi_n_2169), .y(csa_tree_add_14_36_groupi_n_1856));
nor2 csa_tree_add_14_36_groupi_g51002__5266 (.a(csa_tree_add_14_36_groupi_n_1835), .b(csa_tree_add_14_36_groupi_n_1841), .y(csa_tree_add_14_36_groupi_n_1855));
nand2 csa_tree_add_14_36_groupi_g51003__2250 (.a(csa_tree_add_14_36_groupi_n_1777), .b(csa_tree_add_14_36_groupi_n_1843), .y(csa_tree_add_14_36_groupi_n_1854));
nor2 csa_tree_add_14_36_groupi_g51004__6083 (.a(csa_tree_add_14_36_groupi_n_1823), .b(csa_tree_add_14_36_groupi_n_1751), .y(csa_tree_add_14_36_groupi_n_1863));
nand2 csa_tree_add_14_36_groupi_g51006__2703 (.a(csa_tree_add_14_36_groupi_n_1823), .b(csa_tree_add_14_36_groupi_n_1751), .y(csa_tree_add_14_36_groupi_n_2412));
nor2 csa_tree_add_14_36_groupi_g51007__5795 (.a(csa_tree_add_14_36_groupi_n_1832), .b(csa_tree_add_14_36_groupi_n_2174), .y(csa_tree_add_14_36_groupi_n_1861));
nand2 csa_tree_add_14_36_groupi_g51009__7344 (.a(csa_tree_add_14_36_groupi_n_1772), .b(csa_tree_add_14_36_groupi_n_1836), .y(csa_tree_add_14_36_groupi_n_1860));
nand2 csa_tree_add_14_36_groupi_g51010__1840 (.a(csa_tree_add_14_36_groupi_n_1813), .b(csa_tree_add_14_36_groupi_n_1808), .y(csa_tree_add_14_36_groupi_n_1859));
inv csa_tree_add_14_36_groupi_g51013 (.a(csa_tree_add_14_36_groupi_n_1850), .y(csa_tree_add_14_36_groupi_n_2263));
inv csa_tree_add_14_36_groupi_g51014 (.a(csa_tree_add_14_36_groupi_n_2265), .y(csa_tree_add_14_36_groupi_n_1849));
nand2 csa_tree_add_14_36_groupi_g51015__5019 (.a(csa_tree_add_14_36_groupi_n_1822), .b(csa_tree_add_14_36_groupi_n_1819), .y(csa_tree_add_14_36_groupi_n_1848));
nand2 csa_tree_add_14_36_groupi_g51016__1857 (.a(csa_tree_add_14_36_groupi_n_1817), .b(csa_tree_add_14_36_groupi_n_1839), .y(csa_tree_add_14_36_groupi_n_1847));
nand2 csa_tree_add_14_36_groupi_g51017__9906 (.a(n_2683), .b(csa_tree_add_14_36_groupi_n_2214), .y(csa_tree_add_14_36_groupi_n_1846));
nor2 csa_tree_add_14_36_groupi_g51018__8780 (.a(csa_tree_add_14_36_groupi_n_1771), .b(csa_tree_add_14_36_groupi_n_1840), .y(csa_tree_add_14_36_groupi_n_1845));
xor2 csa_tree_add_14_36_groupi_g51019__4296 (.a(csa_tree_add_14_36_groupi_n_1781), .b(csa_tree_add_14_36_groupi_n_1722), .y(csa_tree_add_14_36_groupi_n_2293));
nand2 csa_tree_add_14_36_groupi_g51020__3772 (.a(csa_tree_add_14_36_groupi_n_1824), .b(csa_tree_add_14_36_groupi_n_1756), .y(csa_tree_add_14_36_groupi_n_2410));
xor2 csa_tree_add_14_36_groupi_g51021__1474 (.a(csa_tree_add_14_36_groupi_n_1785), .b(csa_tree_add_14_36_groupi_n_2181), .y(csa_tree_add_14_36_groupi_n_1853));
xor2 csa_tree_add_14_36_groupi_g51024__9682 (.a(csa_tree_add_14_36_groupi_n_1780), .b(csa_tree_add_14_36_groupi_n_2192), .y(csa_tree_add_14_36_groupi_n_1851));
xor2 csa_tree_add_14_36_groupi_g51025__2683 (.a(csa_tree_add_14_36_groupi_n_2209), .b(csa_tree_add_14_36_groupi_n_2213), .y(csa_tree_add_14_36_groupi_n_1844));
nor2 csa_tree_add_14_36_groupi_g51026__1309 (.a(csa_tree_add_14_36_groupi_n_1825), .b(csa_tree_add_14_36_groupi_n_1753), .y(csa_tree_add_14_36_groupi_n_1850));
nand2 csa_tree_add_14_36_groupi_g51027__6877 (.a(csa_tree_add_14_36_groupi_n_1825), .b(csa_tree_add_14_36_groupi_n_1753), .y(csa_tree_add_14_36_groupi_n_2265));
inv csa_tree_add_14_36_groupi_g51028 (.a(csa_tree_add_14_36_groupi_n_1831), .y(csa_tree_add_14_36_groupi_n_1843));
inv csa_tree_add_14_36_groupi_g51029 (.a(csa_tree_add_14_36_groupi_n_1841), .y(csa_tree_add_14_36_groupi_n_1842));
inv csa_tree_add_14_36_groupi_g51030 (.a(csa_tree_add_14_36_groupi_n_1839), .y(csa_tree_add_14_36_groupi_n_1840));
inv csa_tree_add_14_36_groupi_g51031 (.a(csa_tree_add_14_36_groupi_n_1836), .y(csa_tree_add_14_36_groupi_n_1835));
nand2 csa_tree_add_14_36_groupi_g51032__2900 (.a(csa_tree_add_14_36_groupi_n_2209), .b(csa_tree_add_14_36_groupi_n_2213), .y(csa_tree_add_14_36_groupi_n_1834));
nor2 csa_tree_add_14_36_groupi_g51033__2391 (.a(csa_tree_add_14_36_groupi_n_1798), .b(csa_tree_add_14_36_groupi_n_1794), .y(csa_tree_add_14_36_groupi_n_1833));
nor2 csa_tree_add_14_36_groupi_g51034__7675 (.a(csa_tree_add_14_36_groupi_n_2168), .b(csa_tree_add_14_36_groupi_n_2171), .y(csa_tree_add_14_36_groupi_n_1832));
nor2 csa_tree_add_14_36_groupi_g51035__7118 (.a(csa_tree_add_14_36_groupi_n_2209), .b(csa_tree_add_14_36_groupi_n_2213), .y(csa_tree_add_14_36_groupi_n_1831));
nand2 csa_tree_add_14_36_groupi_g51037__8757 (.a(csa_tree_add_14_36_groupi_n_2242), .b(csa_tree_add_14_36_groupi_n_2248), .y(csa_tree_add_14_36_groupi_n_1830));
nor2 csa_tree_add_14_36_groupi_g51038__1786 (.a(csa_tree_add_14_36_groupi_n_1795), .b(csa_tree_add_14_36_groupi_n_1707), .y(csa_tree_add_14_36_groupi_n_1841));
nor2 csa_tree_add_14_36_groupi_g51039__5953 (.a(csa_tree_add_14_36_groupi_n_2169), .b(csa_tree_add_14_36_groupi_n_2171), .y(csa_tree_add_14_36_groupi_n_1839));
nand2 csa_tree_add_14_36_groupi_g51040__5703 (.a(csa_tree_add_14_36_groupi_n_2242), .b(csa_tree_add_14_36_groupi_n_2247), .y(csa_tree_add_14_36_groupi_n_1838));
nor2 csa_tree_add_14_36_groupi_g51041__7114 (.a(csa_tree_add_14_36_groupi_n_2174), .b(csa_tree_add_14_36_groupi_n_2171), .y(csa_tree_add_14_36_groupi_n_1829));
nand2 csa_tree_add_14_36_groupi_g51042__5266 (.a(csa_tree_add_14_36_groupi_n_1804), .b(csa_tree_add_14_36_groupi_n_2165), .y(csa_tree_add_14_36_groupi_n_1828));
nand2 csa_tree_add_14_36_groupi_g51043__2250 (.a(csa_tree_add_14_36_groupi_n_1800), .b(csa_tree_add_14_36_groupi_n_1761), .y(csa_tree_add_14_36_groupi_n_1837));
nand2 csa_tree_add_14_36_groupi_g51044__6083 (.a(csa_tree_add_14_36_groupi_n_2310), .b(csa_tree_add_14_36_groupi_n_2239), .y(csa_tree_add_14_36_groupi_n_1827));
nand2 csa_tree_add_14_36_groupi_g51045__2703 (.a(csa_tree_add_14_36_groupi_n_1795), .b(csa_tree_add_14_36_groupi_n_1707), .y(csa_tree_add_14_36_groupi_n_1836));
inv csa_tree_add_14_36_groupi_g51048 (.a(csa_tree_add_14_36_groupi_n_1821), .y(csa_tree_add_14_36_groupi_n_1822));
inv csa_tree_add_14_36_groupi_g51049 (.a(csa_tree_add_14_36_groupi_n_1819), .y(csa_tree_add_14_36_groupi_n_1820));
inv csa_tree_add_14_36_groupi_g51050 (.a(csa_tree_add_14_36_groupi_n_1818), .y(csa_tree_add_14_36_groupi_n_1817));
nand2 csa_tree_add_14_36_groupi_g51051__5795 (.a(csa_tree_add_14_36_groupi_n_1806), .b(csa_tree_add_14_36_groupi_n_2247), .y(csa_tree_add_14_36_groupi_n_1816));
nor2 csa_tree_add_14_36_groupi_g51052__7344 (.a(csa_tree_add_14_36_groupi_n_1797), .b(csa_tree_add_14_36_groupi_n_1791), .y(csa_tree_add_14_36_groupi_n_1815));
nor2 csa_tree_add_14_36_groupi_g51053__1840 (.a(csa_tree_add_14_36_groupi_n_1806), .b(csa_tree_add_14_36_groupi_n_2247), .y(csa_tree_add_14_36_groupi_n_1814));
nand2 csa_tree_add_14_36_groupi_g51054__5019 (.a(csa_tree_add_14_36_groupi_n_1690), .b(csa_tree_add_14_36_groupi_n_1810), .y(csa_tree_add_14_36_groupi_n_1813));
xor2 csa_tree_add_14_36_groupi_g51055__1857 (.a(csa_tree_add_14_36_groupi_n_1703), .b(csa_tree_add_14_36_groupi_n_1769), .y(result_0__6_));
nand2 csa_tree_add_14_36_groupi_g51056__9906 (.a(csa_tree_add_14_36_groupi_n_1803), .b(csa_tree_add_14_36_groupi_n_1762), .y(csa_tree_add_14_36_groupi_n_1826));
nand2 csa_tree_add_14_36_groupi_g51057__8780 (.a(csa_tree_add_14_36_groupi_n_2247), .b(csa_tree_add_14_36_groupi_n_1807), .y(csa_tree_add_14_36_groupi_n_1812));
xor2 csa_tree_add_14_36_groupi_g51058__4296 (.a(csa_tree_add_14_36_groupi_n_1749), .b(csa_tree_add_14_36_groupi_n_1741), .y(csa_tree_add_14_36_groupi_n_1825));
nand2 csa_tree_add_14_36_groupi_g51059__3772 (.a(csa_tree_add_14_36_groupi_n_1801), .b(csa_tree_add_14_36_groupi_n_1779), .y(csa_tree_add_14_36_groupi_n_1824));
nand2 csa_tree_add_14_36_groupi_g51060__1474 (.a(csa_tree_add_14_36_groupi_n_1788), .b(n_2492), .y(csa_tree_add_14_36_groupi_n_1823));
nor2 csa_tree_add_14_36_groupi_g51061__4547 (.a(csa_tree_add_14_36_groupi_n_1809), .b(csa_tree_add_14_36_groupi_n_1757), .y(csa_tree_add_14_36_groupi_n_1821));
nand2 csa_tree_add_14_36_groupi_g51063__9682 (.a(csa_tree_add_14_36_groupi_n_1787), .b(csa_tree_add_14_36_groupi_n_1727), .y(csa_tree_add_14_36_groupi_n_2294));
nand2 csa_tree_add_14_36_groupi_g51064__2683 (.a(csa_tree_add_14_36_groupi_n_1809), .b(csa_tree_add_14_36_groupi_n_1757), .y(csa_tree_add_14_36_groupi_n_1819));
nor2 csa_tree_add_14_36_groupi_g51065__1309 (.a(csa_tree_add_14_36_groupi_n_1789), .b(csa_tree_add_14_36_groupi_n_1712), .y(csa_tree_add_14_36_groupi_n_1818));
inv csa_tree_add_14_36_groupi_g51069 (.a(csa_tree_add_14_36_groupi_n_2248), .y(csa_tree_add_14_36_groupi_n_1807));
inv csa_tree_add_14_36_groupi_g51070 (.a(csa_tree_add_14_36_groupi_n_1806), .y(csa_tree_add_14_36_groupi_n_1805));
nand2 csa_tree_add_14_36_groupi_g51071__6877 (.a(csa_tree_add_14_36_groupi_n_1769), .b(csa_tree_add_14_36_groupi_n_2163), .y(csa_tree_add_14_36_groupi_n_1804));
nand2 csa_tree_add_14_36_groupi_g51072__2900 (.a(csa_tree_add_14_36_groupi_n_1748), .b(csa_tree_add_14_36_groupi_n_1723), .y(csa_tree_add_14_36_groupi_n_1803));
nand2 csa_tree_add_14_36_groupi_g51073__2391 (.a(csa_tree_add_14_36_groupi_n_1747), .b(csa_tree_add_14_36_groupi_n_1734), .y(csa_tree_add_14_36_groupi_n_1802));
nand2 csa_tree_add_14_36_groupi_g51074__7675 (.a(csa_tree_add_14_36_groupi_n_1764), .b(csa_tree_add_14_36_groupi_n_2192), .y(csa_tree_add_14_36_groupi_n_1801));
nand2 csa_tree_add_14_36_groupi_g51075__7118 (.a(csa_tree_add_14_36_groupi_n_1760), .b(csa_tree_add_14_36_groupi_n_2181), .y(csa_tree_add_14_36_groupi_n_1800));
nor2 csa_tree_add_14_36_groupi_g51077__8757 (.a(csa_tree_add_14_36_groupi_n_1765), .b(n_2476), .y(csa_tree_add_14_36_groupi_n_1811));
nand2 csa_tree_add_14_36_groupi_g51078__1786 (.a(csa_tree_add_14_36_groupi_n_1726), .b(csa_tree_add_14_36_groupi_n_2203), .y(csa_tree_add_14_36_groupi_n_1810));
nand2 csa_tree_add_14_36_groupi_g51079__5953 (.a(csa_tree_add_14_36_groupi_n_1746), .b(csa_tree_add_14_36_groupi_n_1716), .y(csa_tree_add_14_36_groupi_n_1809));
nand2 csa_tree_add_14_36_groupi_g51081__5703 (.a(csa_tree_add_14_36_groupi_n_1725), .b(csa_tree_add_14_36_groupi_n_1778), .y(csa_tree_add_14_36_groupi_n_1808));
nand2 csa_tree_add_14_36_groupi_g51086__7114 (.a(csa_tree_add_14_36_groupi_n_2242), .b(csa_tree_add_14_36_groupi_n_2243), .y(csa_tree_add_14_36_groupi_n_1806));
inv csa_tree_add_14_36_groupi_g51087 (.a(csa_tree_add_14_36_groupi_n_1798), .y(csa_tree_add_14_36_groupi_n_1799));
inv csa_tree_add_14_36_groupi_g51088 (.a(csa_tree_add_14_36_groupi_n_1796), .y(csa_tree_add_14_36_groupi_n_1797));
inv csa_tree_add_14_36_groupi_g51089 (.a(csa_tree_add_14_36_groupi_n_1793), .y(csa_tree_add_14_36_groupi_n_1794));
inv csa_tree_add_14_36_groupi_g51090 (.a(csa_tree_add_14_36_groupi_n_1791), .y(csa_tree_add_14_36_groupi_n_1792));
nor2 csa_tree_add_14_36_groupi_g51091__5266 (.a(csa_tree_add_14_36_groupi_n_1763), .b(csa_tree_add_14_36_groupi_n_1711), .y(csa_tree_add_14_36_groupi_n_1790));
nor2 csa_tree_add_14_36_groupi_g51092__2250 (.a(csa_tree_add_14_36_groupi_n_1699), .b(csa_tree_add_14_36_groupi_n_1768), .y(csa_tree_add_14_36_groupi_n_1789));
nand2 csa_tree_add_14_36_groupi_g51093__6083 (.a(n_2490), .b(csa_tree_add_14_36_groupi_n_2222), .y(csa_tree_add_14_36_groupi_n_1788));
nand2 csa_tree_add_14_36_groupi_g51094__2703 (.a(csa_tree_add_14_36_groupi_n_1749), .b(csa_tree_add_14_36_groupi_n_1724), .y(csa_tree_add_14_36_groupi_n_1787));
nor2 csa_tree_add_14_36_groupi_g51095__5795 (.a(csa_tree_add_14_36_groupi_n_1754), .b(csa_tree_add_14_36_groupi_n_1705), .y(csa_tree_add_14_36_groupi_n_1798));
nor2 csa_tree_add_14_36_groupi_g51096__7344 (.a(csa_tree_add_14_36_groupi_n_1774), .b(csa_tree_add_14_36_groupi_n_1771), .y(csa_tree_add_14_36_groupi_n_1786));
xor2 csa_tree_add_14_36_groupi_g51097__1840 (.a(csa_tree_add_14_36_groupi_n_2184), .b(csa_tree_add_14_36_groupi_n_2191), .y(csa_tree_add_14_36_groupi_n_1785));
nand2 csa_tree_add_14_36_groupi_g51098__5019 (.a(csa_tree_add_14_36_groupi_n_1758), .b(csa_tree_add_14_36_groupi_n_2236), .y(csa_tree_add_14_36_groupi_n_1796));
nand2 csa_tree_add_14_36_groupi_g51101__8780 (.a(csa_tree_add_14_36_groupi_n_1776), .b(csa_tree_add_14_36_groupi_n_1772), .y(csa_tree_add_14_36_groupi_n_1782));
xor2 csa_tree_add_14_36_groupi_g51102__4296 (.a(csa_tree_add_14_36_groupi_n_1721), .b(csa_tree_add_14_36_groupi_n_2205), .y(csa_tree_add_14_36_groupi_n_1781));
xor2 csa_tree_add_14_36_groupi_g51104__1474 (.a(csa_tree_add_14_36_groupi_n_1710), .b(csa_tree_add_14_36_groupi_n_2179), .y(csa_tree_add_14_36_groupi_n_1795));
xor2 csa_tree_add_14_36_groupi_g51105__4547 (.a(csa_tree_add_14_36_groupi_n_2196), .b(csa_tree_add_14_36_groupi_n_2186), .y(csa_tree_add_14_36_groupi_n_1780));
nand2 csa_tree_add_14_36_groupi_g51106__9682 (.a(csa_tree_add_14_36_groupi_n_1754), .b(csa_tree_add_14_36_groupi_n_1705), .y(csa_tree_add_14_36_groupi_n_1793));
nor2 csa_tree_add_14_36_groupi_g51107__2683 (.a(csa_tree_add_14_36_groupi_n_1758), .b(csa_tree_add_14_36_groupi_n_2236), .y(csa_tree_add_14_36_groupi_n_1791));
inv csa_tree_add_14_36_groupi_g51108 (.a(csa_tree_add_14_36_groupi_n_1766), .y(csa_tree_add_14_36_groupi_n_1779));
inv csa_tree_add_14_36_groupi_g51109 (.a(csa_tree_add_14_36_groupi_n_2203), .y(csa_tree_add_14_36_groupi_n_1778));
inv csa_tree_add_14_36_groupi_g51110 (.a(csa_tree_add_14_36_groupi_n_1775), .y(csa_tree_add_14_36_groupi_n_1776));
inv csa_tree_add_14_36_groupi_g51111 (.a(csa_tree_add_14_36_groupi_n_1773), .y(csa_tree_add_14_36_groupi_n_1774));
inv csa_tree_add_14_36_groupi_g51112 (.a(csa_tree_add_14_36_groupi_n_1771), .y(csa_tree_add_14_36_groupi_n_1770));
inv csa_tree_add_14_36_groupi_g51113 (.a(csa_tree_add_14_36_groupi_n_1769), .y(csa_tree_add_14_36_groupi_n_1768));
nor2 csa_tree_add_14_36_groupi_g51114__1309 (.a(csa_tree_add_14_36_groupi_n_1569), .b(csa_tree_add_14_36_groupi_n_1728), .y(csa_tree_add_14_36_groupi_n_1767));
nor2 csa_tree_add_14_36_groupi_g51115__6877 (.a(csa_tree_add_14_36_groupi_n_2196), .b(csa_tree_add_14_36_groupi_n_2186), .y(csa_tree_add_14_36_groupi_n_1766));
nor2 csa_tree_add_14_36_groupi_g51116__2900 (.a(n_2478), .b(csa_tree_add_14_36_groupi_n_2218), .y(csa_tree_add_14_36_groupi_n_1765));
nand2 csa_tree_add_14_36_groupi_g51117__2391 (.a(csa_tree_add_14_36_groupi_n_2196), .b(csa_tree_add_14_36_groupi_n_2186), .y(csa_tree_add_14_36_groupi_n_1764));
nor2 csa_tree_add_14_36_groupi_g51118__7675 (.a(csa_tree_add_14_36_groupi_n_1735), .b(csa_tree_add_14_36_groupi_n_130), .y(csa_tree_add_14_36_groupi_n_1763));
nand2 csa_tree_add_14_36_groupi_g51120__7118 (.a(csa_tree_add_14_36_groupi_n_1721), .b(csa_tree_add_14_36_groupi_n_1701), .y(csa_tree_add_14_36_groupi_n_1762));
nand2 csa_tree_add_14_36_groupi_g51122__8757 (.a(csa_tree_add_14_36_groupi_n_1627), .b(csa_tree_add_14_36_groupi_n_2191), .y(csa_tree_add_14_36_groupi_n_1761));
nand2 csa_tree_add_14_36_groupi_g51125__1786 (.a(csa_tree_add_14_36_groupi_n_2184), .b(csa_tree_add_14_36_groupi_n_1737), .y(csa_tree_add_14_36_groupi_n_1760));
nand2 csa_tree_add_14_36_groupi_g51126__5953 (.a(csa_tree_add_14_36_groupi_n_1719), .b(csa_tree_add_14_36_groupi_n_1697), .y(csa_tree_add_14_36_groupi_n_1777));
nor2 csa_tree_add_14_36_groupi_g51127__5703 (.a(csa_tree_add_14_36_groupi_n_1729), .b(csa_tree_add_14_36_groupi_n_2320), .y(csa_tree_add_14_36_groupi_n_1775));
nand2 csa_tree_add_14_36_groupi_g51128__7114 (.a(csa_tree_add_14_36_groupi_n_2321), .b(csa_tree_add_14_36_groupi_n_2173), .y(csa_tree_add_14_36_groupi_n_1773));
nand2 csa_tree_add_14_36_groupi_g51129__5266 (.a(csa_tree_add_14_36_groupi_n_1729), .b(csa_tree_add_14_36_groupi_n_2320), .y(csa_tree_add_14_36_groupi_n_1772));
nor2 csa_tree_add_14_36_groupi_g51131__2250 (.a(csa_tree_add_14_36_groupi_n_2321), .b(csa_tree_add_14_36_groupi_n_2173), .y(csa_tree_add_14_36_groupi_n_1771));
nand2 csa_tree_add_14_36_groupi_g51132__6083 (.a(csa_tree_add_14_36_groupi_n_2160), .b(csa_tree_add_14_36_groupi_n_2162), .y(csa_tree_add_14_36_groupi_n_1769));
nand2 csa_tree_add_14_36_groupi_g51134__2703 (.a(csa_tree_add_14_36_groupi_n_1720), .b(csa_tree_add_14_36_groupi_n_2205), .y(csa_tree_add_14_36_groupi_n_1748));
nand2 csa_tree_add_14_36_groupi_g51135__5795 (.a(csa_tree_add_14_36_groupi_n_1740), .b(csa_tree_add_14_36_groupi_n_1497), .y(csa_tree_add_14_36_groupi_n_1747));
nand2 csa_tree_add_14_36_groupi_g51136__7344 (.a(csa_tree_add_14_36_groupi_n_1718), .b(csa_tree_add_14_36_groupi_n_2314), .y(csa_tree_add_14_36_groupi_n_1746));
nand2 csa_tree_add_14_36_groupi_g51138__5019 (.a(n_2486), .b(csa_tree_add_14_36_groupi_n_2249), .y(csa_tree_add_14_36_groupi_n_1744));
nand2 csa_tree_add_14_36_groupi_g51139__1857 (.a(csa_tree_add_14_36_groupi_n_1691), .b(csa_tree_add_14_36_groupi_n_2261), .y(csa_tree_add_14_36_groupi_n_1743));
xor2 csa_tree_add_14_36_groupi_g51140__9906 (.a(csa_tree_add_14_36_groupi_n_1661), .b(csa_tree_add_14_36_groupi_n_2161), .y(result_0__5_));
xor2 csa_tree_add_14_36_groupi_g51141__8780 (.a(n_2551), .b(csa_tree_add_14_36_groupi_n_1582), .y(csa_tree_add_14_36_groupi_n_1742));
nor2 csa_tree_add_14_36_groupi_g51143__3772 (.a(csa_tree_add_14_36_groupi_n_1731), .b(csa_tree_add_14_36_groupi_n_1612), .y(csa_tree_add_14_36_groupi_n_1758));
nand2 csa_tree_add_14_36_groupi_g51144__1474 (.a(csa_tree_add_14_36_groupi_n_1727), .b(csa_tree_add_14_36_groupi_n_1724), .y(csa_tree_add_14_36_groupi_n_1741));
xor2 csa_tree_add_14_36_groupi_g51145__4547 (.a(csa_tree_add_14_36_groupi_n_1637), .b(csa_tree_add_14_36_groupi_n_2229), .y(csa_tree_add_14_36_groupi_n_1757));
xor2 csa_tree_add_14_36_groupi_g51146__9682 (.a(n_2468), .b(csa_tree_add_14_36_groupi_n_2189), .y(csa_tree_add_14_36_groupi_n_1756));
xor2 csa_tree_add_14_36_groupi_g51148__1309 (.a(csa_tree_add_14_36_groupi_n_1673), .b(csa_tree_add_14_36_groupi_n_2170), .y(csa_tree_add_14_36_groupi_n_1754));
nand2 csa_tree_add_14_36_groupi_g51149__6877 (.a(csa_tree_add_14_36_groupi_n_1713), .b(n_2470), .y(csa_tree_add_14_36_groupi_n_1753));
xor2 csa_tree_add_14_36_groupi_g51151__2391 (.a(csa_tree_add_14_36_groupi_n_1674), .b(csa_tree_add_14_36_groupi_n_2224), .y(csa_tree_add_14_36_groupi_n_1751));
xor2 csa_tree_add_14_36_groupi_g51153__7118 (.a(csa_tree_add_14_36_groupi_n_1676), .b(csa_tree_add_14_36_groupi_n_2193), .y(csa_tree_add_14_36_groupi_n_1749));
inv csa_tree_add_14_36_groupi_g51154 (.a(n_2550), .y(csa_tree_add_14_36_groupi_n_1740));
inv csa_tree_add_14_36_groupi_g51156 (.a(csa_tree_add_14_36_groupi_n_2191), .y(csa_tree_add_14_36_groupi_n_1737));
nand2 csa_tree_add_14_36_groupi_g51158__8757 (.a(n_2551), .b(n_2547), .y(csa_tree_add_14_36_groupi_n_1734));
nand2 csa_tree_add_14_36_groupi_g51160__1786 (.a(csa_tree_add_14_36_groupi_n_1708), .b(csa_tree_add_14_36_groupi_n_2241), .y(csa_tree_add_14_36_groupi_n_1733));
nor2 csa_tree_add_14_36_groupi_g51162__5703 (.a(csa_tree_add_14_36_groupi_n_1611), .b(csa_tree_add_14_36_groupi_n_2229), .y(csa_tree_add_14_36_groupi_n_1731));
nand2 csa_tree_add_14_36_groupi_g51166__7114 (.a(csa_tree_add_14_36_groupi_n_2237), .b(csa_tree_add_14_36_groupi_n_2232), .y(csa_tree_add_14_36_groupi_n_2261));
nor2 csa_tree_add_14_36_groupi_g51167__5266 (.a(csa_tree_add_14_36_groupi_n_2250), .b(csa_tree_add_14_36_groupi_n_2245), .y(csa_tree_add_14_36_groupi_n_1730));
nor2 csa_tree_add_14_36_groupi_g51168__2250 (.a(csa_tree_add_14_36_groupi_n_1662), .b(csa_tree_add_14_36_groupi_n_1696), .y(csa_tree_add_14_36_groupi_n_1738));
nand2 csa_tree_add_14_36_groupi_g51171__6083 (.a(csa_tree_add_14_36_groupi_n_2240), .b(csa_tree_add_14_36_groupi_n_1702), .y(csa_tree_add_14_36_groupi_n_1735));
inv csa_tree_add_14_36_groupi_g51176 (.a(csa_tree_add_14_36_groupi_n_1725), .y(csa_tree_add_14_36_groupi_n_1726));
inv csa_tree_add_14_36_groupi_g51177 (.a(csa_tree_add_14_36_groupi_n_1722), .y(csa_tree_add_14_36_groupi_n_1723));
inv csa_tree_add_14_36_groupi_g51178 (.a(csa_tree_add_14_36_groupi_n_1721), .y(csa_tree_add_14_36_groupi_n_1720));
nand2 csa_tree_add_14_36_groupi_g51179__2703 (.a(csa_tree_add_14_36_groupi_n_1709), .b(csa_tree_add_14_36_groupi_n_2207), .y(csa_tree_add_14_36_groupi_n_1719));
nand2 csa_tree_add_14_36_groupi_g51180__5795 (.a(csa_tree_add_14_36_groupi_n_1624), .b(csa_tree_add_14_36_groupi_n_2224), .y(csa_tree_add_14_36_groupi_n_1718));
nand2 csa_tree_add_14_36_groupi_g51181__7344 (.a(csa_tree_add_14_36_groupi_n_2244), .b(csa_tree_add_14_36_groupi_n_1672), .y(csa_tree_add_14_36_groupi_n_1717));
nand2 csa_tree_add_14_36_groupi_g51182__1840 (.a(csa_tree_add_14_36_groupi_n_2226), .b(csa_tree_add_14_36_groupi_n_1700), .y(csa_tree_add_14_36_groupi_n_1716));
xor2 csa_tree_add_14_36_groupi_g51183__5019 (.a(n_2543), .b(csa_tree_add_14_36_groupi_n_1600), .y(csa_tree_add_14_36_groupi_n_1715));
xor2 csa_tree_add_14_36_groupi_g51184__1857 (.a(csa_tree_add_14_36_groupi_n_1472), .b(csa_tree_add_14_36_groupi_n_1643), .y(csa_tree_add_14_36_groupi_n_1714));
nand2 csa_tree_add_14_36_groupi_g51185__9906 (.a(n_2472), .b(csa_tree_add_14_36_groupi_n_2189), .y(csa_tree_add_14_36_groupi_n_1713));
nand2 csa_tree_add_14_36_groupi_g51186__8780 (.a(csa_tree_add_14_36_groupi_n_1680), .b(csa_tree_add_14_36_groupi_n_2164), .y(csa_tree_add_14_36_groupi_n_1712));
nor2 csa_tree_add_14_36_groupi_g51187__4296 (.a(csa_tree_add_14_36_groupi_n_2240), .b(csa_tree_add_14_36_groupi_n_1702), .y(csa_tree_add_14_36_groupi_n_1711));
nand2 csa_tree_add_14_36_groupi_g51188__3772 (.a(csa_tree_add_14_36_groupi_n_1681), .b(csa_tree_add_14_36_groupi_n_1647), .y(csa_tree_add_14_36_groupi_n_1729));
xor2 csa_tree_add_14_36_groupi_g51189__1474 (.a(csa_tree_add_14_36_groupi_n_1640), .b(csa_tree_add_14_36_groupi_n_1403), .y(csa_tree_add_14_36_groupi_n_1728));
nand2 csa_tree_add_14_36_groupi_g51190__4547 (.a(csa_tree_add_14_36_groupi_n_1629), .b(csa_tree_add_14_36_groupi_n_2200), .y(csa_tree_add_14_36_groupi_n_1727));
xor2 csa_tree_add_14_36_groupi_g51191__9682 (.a(csa_tree_add_14_36_groupi_n_1645), .b(csa_tree_add_14_36_groupi_n_2204), .y(csa_tree_add_14_36_groupi_n_1725));
nand2 csa_tree_add_14_36_groupi_g51192__2683 (.a(csa_tree_add_14_36_groupi_n_2202), .b(csa_tree_add_14_36_groupi_n_1706), .y(csa_tree_add_14_36_groupi_n_1724));
xor2 csa_tree_add_14_36_groupi_g51193__1309 (.a(csa_tree_add_14_36_groupi_n_2319), .b(csa_tree_add_14_36_groupi_n_2182), .y(csa_tree_add_14_36_groupi_n_1710));
nor2 csa_tree_add_14_36_groupi_g51194__6877 (.a(csa_tree_add_14_36_groupi_n_1682), .b(csa_tree_add_14_36_groupi_n_1644), .y(csa_tree_add_14_36_groupi_n_1722));
xor2 csa_tree_add_14_36_groupi_g51195__2900 (.a(csa_tree_add_14_36_groupi_n_1642), .b(csa_tree_add_14_36_groupi_n_2201), .y(csa_tree_add_14_36_groupi_n_1721));
inv csa_tree_add_14_36_groupi_g51196 (.a(csa_tree_add_14_36_groupi_n_1698), .y(csa_tree_add_14_36_groupi_n_1709));
inv csa_tree_add_14_36_groupi_g51197 (.a(csa_tree_add_14_36_groupi_n_2244), .y(csa_tree_add_14_36_groupi_n_1708));
inv csa_tree_add_14_36_groupi_g51198 (.a(csa_tree_add_14_36_groupi_n_2200), .y(csa_tree_add_14_36_groupi_n_1706));
inv csa_tree_add_14_36_groupi_g51199 (.a(csa_tree_add_14_36_groupi_n_1695), .y(csa_tree_add_14_36_groupi_n_1704));
inv csa_tree_add_14_36_groupi_g51200 (.a(csa_tree_add_14_36_groupi_n_1694), .y(csa_tree_add_14_36_groupi_n_1703));
inv csa_tree_add_14_36_groupi_g51201 (.a(csa_tree_add_14_36_groupi_n_2245), .y(csa_tree_add_14_36_groupi_n_1702));
inv csa_tree_add_14_36_groupi_g51202 (.a(csa_tree_add_14_36_groupi_n_2205), .y(csa_tree_add_14_36_groupi_n_1701));
inv csa_tree_add_14_36_groupi_g51203 (.a(csa_tree_add_14_36_groupi_n_2224), .y(csa_tree_add_14_36_groupi_n_1700));
nand2 csa_tree_add_14_36_groupi_g51204__2391 (.a(csa_tree_add_14_36_groupi_n_2303), .b(csa_tree_add_14_36_groupi_n_2163), .y(csa_tree_add_14_36_groupi_n_1699));
nor2 csa_tree_add_14_36_groupi_g51205__7675 (.a(csa_tree_add_14_36_groupi_n_2216), .b(csa_tree_add_14_36_groupi_n_2204), .y(csa_tree_add_14_36_groupi_n_1698));
nand2 csa_tree_add_14_36_groupi_g51206__7118 (.a(csa_tree_add_14_36_groupi_n_2216), .b(csa_tree_add_14_36_groupi_n_2204), .y(csa_tree_add_14_36_groupi_n_1697));
nor2 csa_tree_add_14_36_groupi_g51209__8757 (.a(csa_tree_add_14_36_groupi_n_2185), .b(csa_tree_add_14_36_groupi_n_2182), .y(csa_tree_add_14_36_groupi_n_1696));
nor2 csa_tree_add_14_36_groupi_g51211__1786 (.a(csa_tree_add_14_36_groupi_n_2183), .b(csa_tree_add_14_36_groupi_n_2180), .y(csa_tree_add_14_36_groupi_n_1707));
nor2 csa_tree_add_14_36_groupi_g51213__5953 (.a(csa_tree_add_14_36_groupi_n_2175), .b(csa_tree_add_14_36_groupi_n_2172), .y(csa_tree_add_14_36_groupi_n_1705));
nand2 csa_tree_add_14_36_groupi_g51215__5703 (.a(csa_tree_add_14_36_groupi_n_2303), .b(csa_tree_add_14_36_groupi_n_2164), .y(csa_tree_add_14_36_groupi_n_1695));
nand2 csa_tree_add_14_36_groupi_g51216__7114 (.a(csa_tree_add_14_36_groupi_n_2165), .b(csa_tree_add_14_36_groupi_n_2163), .y(csa_tree_add_14_36_groupi_n_1694));
nand2 csa_tree_add_14_36_groupi_g51217__5266 (.a(csa_tree_add_14_36_groupi_n_2168), .b(csa_tree_add_14_36_groupi_n_1671), .y(csa_tree_add_14_36_groupi_n_1693));
inv csa_tree_add_14_36_groupi_g51224 (.a(csa_tree_add_14_36_groupi_n_2266), .y(csa_tree_add_14_36_groupi_n_1691));
nand2 csa_tree_add_14_36_groupi_g51225__2250 (.a(csa_tree_add_14_36_groupi_n_1664), .b(csa_tree_add_14_36_groupi_n_1617), .y(csa_tree_add_14_36_groupi_n_1688));
nor2 csa_tree_add_14_36_groupi_g51226__6083 (.a(csa_tree_add_14_36_groupi_n_1666), .b(csa_tree_add_14_36_groupi_n_1602), .y(csa_tree_add_14_36_groupi_n_1687));
xor2 csa_tree_add_14_36_groupi_g51227__2703 (.a(csa_tree_add_14_36_groupi_n_1496), .b(csa_tree_add_14_36_groupi_n_1577), .y(csa_tree_add_14_36_groupi_n_1686));
nand2 csa_tree_add_14_36_groupi_g51228__5795 (.a(csa_tree_add_14_36_groupi_n_1669), .b(csa_tree_add_14_36_groupi_n_1621), .y(csa_tree_add_14_36_groupi_n_1685));
nand2 csa_tree_add_14_36_groupi_g51229__7344 (.a(csa_tree_add_14_36_groupi_n_1663), .b(csa_tree_add_14_36_groupi_n_1608), .y(csa_tree_add_14_36_groupi_n_1684));
xor2 csa_tree_add_14_36_groupi_g51230__1840 (.a(csa_tree_add_14_36_groupi_n_1543), .b(csa_tree_add_14_36_groupi_n_1580), .y(csa_tree_add_14_36_groupi_n_1683));
nor2 csa_tree_add_14_36_groupi_g51231__5019 (.a(csa_tree_add_14_36_groupi_n_1639), .b(csa_tree_add_14_36_groupi_n_2193), .y(csa_tree_add_14_36_groupi_n_1682));
nand2 csa_tree_add_14_36_groupi_g51232__1857 (.a(csa_tree_add_14_36_groupi_n_1646), .b(csa_tree_add_14_36_groupi_n_2170), .y(csa_tree_add_14_36_groupi_n_1681));
nand2 csa_tree_add_14_36_groupi_g51233__9906 (.a(csa_tree_add_14_36_groupi_n_2303), .b(csa_tree_add_14_36_groupi_n_1670), .y(csa_tree_add_14_36_groupi_n_1680));
xor2 csa_tree_add_14_36_groupi_g51234__8780 (.a(csa_tree_add_14_36_groupi_n_1583), .b(csa_tree_add_14_36_groupi_n_1474), .y(csa_tree_add_14_36_groupi_n_1679));
xor2 csa_tree_add_14_36_groupi_g51235__4296 (.a(csa_tree_add_14_36_groupi_n_1498), .b(csa_tree_add_14_36_groupi_n_1610), .y(csa_tree_add_14_36_groupi_n_1678));
xor2 csa_tree_add_14_36_groupi_g51236__3772 (.a(csa_tree_add_14_36_groupi_n_1578), .b(csa_tree_add_14_36_groupi_n_1512), .y(csa_tree_add_14_36_groupi_n_1677));
xor2 csa_tree_add_14_36_groupi_g51238__4547 (.a(csa_tree_add_14_36_groupi_n_2255), .b(csa_tree_add_14_36_groupi_n_2141), .y(csa_tree_add_14_36_groupi_n_1676));
xor2 csa_tree_add_14_36_groupi_g51240__2683 (.a(csa_tree_add_14_36_groupi_n_2314), .b(csa_tree_add_14_36_groupi_n_2226), .y(csa_tree_add_14_36_groupi_n_1674));
xor2 csa_tree_add_14_36_groupi_g51241__1309 (.a(csa_tree_add_14_36_groupi_n_1524), .b(csa_tree_add_14_36_groupi_n_2178), .y(csa_tree_add_14_36_groupi_n_1673));
xor2 csa_tree_add_14_36_groupi_g51242__6877 (.a(csa_tree_add_14_36_groupi_n_1526), .b(csa_tree_add_14_36_groupi_n_2238), .y(csa_tree_add_14_36_groupi_n_2266));
nor2 csa_tree_add_14_36_groupi_g51243__2900 (.a(csa_tree_add_14_36_groupi_n_1655), .b(csa_tree_add_14_36_groupi_n_1579), .y(csa_tree_add_14_36_groupi_n_1690));
inv csa_tree_add_14_36_groupi_g51245 (.a(csa_tree_add_14_36_groupi_n_2241), .y(csa_tree_add_14_36_groupi_n_1672));
inv csa_tree_add_14_36_groupi_g51246 (.a(csa_tree_add_14_36_groupi_n_2169), .y(csa_tree_add_14_36_groupi_n_1671));
inv csa_tree_add_14_36_groupi_g51247 (.a(csa_tree_add_14_36_groupi_n_2165), .y(csa_tree_add_14_36_groupi_n_1670));
nand2 csa_tree_add_14_36_groupi_g51248__7675 (.a(csa_tree_add_14_36_groupi_n_1635), .b(csa_tree_add_14_36_groupi_n_2286), .y(csa_tree_add_14_36_groupi_n_1669));
nand2 csa_tree_add_14_36_groupi_g51250__7118 (.a(csa_tree_add_14_36_groupi_n_1599), .b(csa_tree_add_14_36_groupi_n_1558), .y(csa_tree_add_14_36_groupi_n_1668));
nand2 csa_tree_add_14_36_groupi_g51252__8757 (.a(csa_tree_add_14_36_groupi_n_1636), .b(csa_tree_add_14_36_groupi_n_1568), .y(csa_tree_add_14_36_groupi_n_1667));
nor2 csa_tree_add_14_36_groupi_g51253__1786 (.a(n_2431), .b(csa_tree_add_14_36_groupi_n_1358), .y(csa_tree_add_14_36_groupi_n_1666));
nand2 csa_tree_add_14_36_groupi_g51256__5703 (.a(csa_tree_add_14_36_groupi_n_1633), .b(csa_tree_add_14_36_groupi_n_1403), .y(csa_tree_add_14_36_groupi_n_1664));
nand2 csa_tree_add_14_36_groupi_g51257__7114 (.a(csa_tree_add_14_36_groupi_n_1597), .b(csa_tree_add_14_36_groupi_n_1494), .y(csa_tree_add_14_36_groupi_n_1663));
nor2 csa_tree_add_14_36_groupi_g51258__5266 (.a(csa_tree_add_14_36_groupi_n_2319), .b(csa_tree_add_14_36_groupi_n_2179), .y(csa_tree_add_14_36_groupi_n_1662));
nor2 csa_tree_add_14_36_groupi_g51261__2250 (.a(csa_tree_add_14_36_groupi_n_2159), .b(csa_tree_add_14_36_groupi_n_2166), .y(csa_tree_add_14_36_groupi_n_1661));
nand2 csa_tree_add_14_36_groupi_g51272__6083 (.a(csa_tree_add_14_36_groupi_n_1609), .b(csa_tree_add_14_36_groupi_n_1559), .y(csa_tree_add_14_36_groupi_n_1657));
nand2 csa_tree_add_14_36_groupi_g51273__2703 (.a(csa_tree_add_14_36_groupi_n_1634), .b(csa_tree_add_14_36_groupi_n_1600), .y(csa_tree_add_14_36_groupi_n_1656));
nor2 csa_tree_add_14_36_groupi_g51274__5795 (.a(csa_tree_add_14_36_groupi_n_1581), .b(csa_tree_add_14_36_groupi_n_2201), .y(csa_tree_add_14_36_groupi_n_1655));
nand2 csa_tree_add_14_36_groupi_g51275__7344 (.a(csa_tree_add_14_36_groupi_n_1482), .b(csa_tree_add_14_36_groupi_n_1625), .y(csa_tree_add_14_36_groupi_n_1654));
nand2 csa_tree_add_14_36_groupi_g51276__1840 (.a(csa_tree_add_14_36_groupi_n_1596), .b(csa_tree_add_14_36_groupi_n_1553), .y(csa_tree_add_14_36_groupi_n_1653));
nand2 csa_tree_add_14_36_groupi_g51277__5019 (.a(csa_tree_add_14_36_groupi_n_1594), .b(csa_tree_add_14_36_groupi_n_1538), .y(csa_tree_add_14_36_groupi_n_1652));
nand2 csa_tree_add_14_36_groupi_g51278__1857 (.a(csa_tree_add_14_36_groupi_n_1472), .b(csa_tree_add_14_36_groupi_n_1604), .y(csa_tree_add_14_36_groupi_n_1651));
nand2 csa_tree_add_14_36_groupi_g51279__9906 (.a(csa_tree_add_14_36_groupi_n_1601), .b(n_2438), .y(csa_tree_add_14_36_groupi_n_1650));
nand2 csa_tree_add_14_36_groupi_g51280__8780 (.a(csa_tree_add_14_36_groupi_n_1588), .b(csa_tree_add_14_36_groupi_n_1551), .y(csa_tree_add_14_36_groupi_n_1649));
xor2 csa_tree_add_14_36_groupi_g51281__4296 (.a(csa_tree_add_14_36_groupi_n_1359), .b(csa_tree_add_14_36_groupi_n_1527), .y(csa_tree_add_14_36_groupi_n_1648));
nand2 csa_tree_add_14_36_groupi_g51284__4547 (.a(csa_tree_add_14_36_groupi_n_1524), .b(csa_tree_add_14_36_groupi_n_2178), .y(csa_tree_add_14_36_groupi_n_1647));
nand2 csa_tree_add_14_36_groupi_g51285__9682 (.a(csa_tree_add_14_36_groupi_n_2176), .b(csa_tree_add_14_36_groupi_n_1631), .y(csa_tree_add_14_36_groupi_n_1646));
xor2 csa_tree_add_14_36_groupi_g51286__2683 (.a(csa_tree_add_14_36_groupi_n_2216), .b(csa_tree_add_14_36_groupi_n_2207), .y(csa_tree_add_14_36_groupi_n_1645));
nor2 csa_tree_add_14_36_groupi_g51287__1309 (.a(csa_tree_add_14_36_groupi_n_2255), .b(csa_tree_add_14_36_groupi_n_1630), .y(csa_tree_add_14_36_groupi_n_1644));
nand2 csa_tree_add_14_36_groupi_g51288__6877 (.a(csa_tree_add_14_36_groupi_n_1605), .b(csa_tree_add_14_36_groupi_n_1604), .y(csa_tree_add_14_36_groupi_n_1643));
xor2 csa_tree_add_14_36_groupi_g51289__2900 (.a(csa_tree_add_14_36_groupi_n_65), .b(csa_tree_add_14_36_groupi_n_2138), .y(csa_tree_add_14_36_groupi_n_1642));
xor2 csa_tree_add_14_36_groupi_g51291__7675 (.a(csa_tree_add_14_36_groupi_n_1542), .b(csa_tree_add_14_36_groupi_n_1251), .y(csa_tree_add_14_36_groupi_n_1640));
nor2 csa_tree_add_14_36_groupi_g51292__7118 (.a(csa_tree_add_14_36_groupi_n_1521), .b(csa_tree_add_14_36_groupi_n_2141), .y(csa_tree_add_14_36_groupi_n_1639));
xor2 csa_tree_add_14_36_groupi_g51294__1786 (.a(csa_tree_add_14_36_groupi_n_87), .b(csa_tree_add_14_36_groupi_n_2223), .y(csa_tree_add_14_36_groupi_n_1637));
inv csa_tree_add_14_36_groupi_g51295 (.a(csa_tree_add_14_36_groupi_n_1622), .y(csa_tree_add_14_36_groupi_n_1636));
inv csa_tree_add_14_36_groupi_g51296 (.a(csa_tree_add_14_36_groupi_n_1620), .y(csa_tree_add_14_36_groupi_n_1635));
inv csa_tree_add_14_36_groupi_g51297 (.a(csa_tree_add_14_36_groupi_n_1618), .y(csa_tree_add_14_36_groupi_n_1634));
inv csa_tree_add_14_36_groupi_g51298 (.a(csa_tree_add_14_36_groupi_n_1616), .y(csa_tree_add_14_36_groupi_n_1633));
inv csa_tree_add_14_36_groupi_g51300 (.a(csa_tree_add_14_36_groupi_n_2178), .y(csa_tree_add_14_36_groupi_n_1631));
inv csa_tree_add_14_36_groupi_g51301 (.a(csa_tree_add_14_36_groupi_n_2141), .y(csa_tree_add_14_36_groupi_n_1630));
inv csa_tree_add_14_36_groupi_g51302 (.a(csa_tree_add_14_36_groupi_n_2202), .y(csa_tree_add_14_36_groupi_n_1629));
inv csa_tree_add_14_36_groupi_g51304 (.a(csa_tree_add_14_36_groupi_n_2184), .y(csa_tree_add_14_36_groupi_n_1627));
inv csa_tree_add_14_36_groupi_g51306 (.a(csa_tree_add_14_36_groupi_n_2238), .y(csa_tree_add_14_36_groupi_n_1625));
inv csa_tree_add_14_36_groupi_g51307 (.a(csa_tree_add_14_36_groupi_n_2226), .y(csa_tree_add_14_36_groupi_n_1624));
nor2 csa_tree_add_14_36_groupi_g51308__5953 (.a(csa_tree_add_14_36_groupi_n_1571), .b(csa_tree_add_14_36_groupi_n_1549), .y(csa_tree_add_14_36_groupi_n_1623));
nor2 csa_tree_add_14_36_groupi_g51311__5703 (.a(csa_tree_add_14_36_groupi_n_1498), .b(csa_tree_add_14_36_groupi_n_1574), .y(csa_tree_add_14_36_groupi_n_1622));
nand2 csa_tree_add_14_36_groupi_g51312__7114 (.a(csa_tree_add_14_36_groupi_n_2288), .b(csa_tree_add_14_36_groupi_n_2287), .y(csa_tree_add_14_36_groupi_n_1621));
nor2 csa_tree_add_14_36_groupi_g51313__5266 (.a(csa_tree_add_14_36_groupi_n_2288), .b(csa_tree_add_14_36_groupi_n_2287), .y(csa_tree_add_14_36_groupi_n_1620));
nand2 csa_tree_add_14_36_groupi_g51314__2250 (.a(n_2544), .b(csa_tree_add_14_36_groupi_n_2064), .y(csa_tree_add_14_36_groupi_n_1619));
nor2 csa_tree_add_14_36_groupi_g51315__6083 (.a(n_2544), .b(csa_tree_add_14_36_groupi_n_2064), .y(csa_tree_add_14_36_groupi_n_1618));
nand2 csa_tree_add_14_36_groupi_g51316__2703 (.a(csa_tree_add_14_36_groupi_n_1542), .b(csa_tree_add_14_36_groupi_n_1251), .y(csa_tree_add_14_36_groupi_n_1617));
nor2 csa_tree_add_14_36_groupi_g51317__5795 (.a(csa_tree_add_14_36_groupi_n_1542), .b(csa_tree_add_14_36_groupi_n_1251), .y(csa_tree_add_14_36_groupi_n_1616));
nor2 csa_tree_add_14_36_groupi_g51318__7344 (.a(csa_tree_add_14_36_groupi_n_1555), .b(n_2624), .y(csa_tree_add_14_36_groupi_n_1615));
nand2 csa_tree_add_14_36_groupi_g51319__1840 (.a(csa_tree_add_14_36_groupi_n_1520), .b(csa_tree_add_14_36_groupi_n_1547), .y(csa_tree_add_14_36_groupi_n_1614));
nand2 csa_tree_add_14_36_groupi_g51320__5019 (.a(csa_tree_add_14_36_groupi_n_1519), .b(csa_tree_add_14_36_groupi_n_1548), .y(csa_tree_add_14_36_groupi_n_1613));
nor2 csa_tree_add_14_36_groupi_g51322__1857 (.a(csa_tree_add_14_36_groupi_n_87), .b(csa_tree_add_14_36_groupi_n_1573), .y(csa_tree_add_14_36_groupi_n_1612));
nor2 csa_tree_add_14_36_groupi_g51324__9906 (.a(csa_tree_add_14_36_groupi_n_2309), .b(csa_tree_add_14_36_groupi_n_2223), .y(csa_tree_add_14_36_groupi_n_1611));
nand2 csa_tree_add_14_36_groupi_g51326__8780 (.a(csa_tree_add_14_36_groupi_n_1575), .b(csa_tree_add_14_36_groupi_n_1568), .y(csa_tree_add_14_36_groupi_n_1610));
inv csa_tree_add_14_36_groupi_g51339 (.a(csa_tree_add_14_36_groupi_n_1598), .y(csa_tree_add_14_36_groupi_n_1609));
inv csa_tree_add_14_36_groupi_g51340 (.a(csa_tree_add_14_36_groupi_n_1595), .y(csa_tree_add_14_36_groupi_n_1608));
inv csa_tree_add_14_36_groupi_g51341 (.a(csa_tree_add_14_36_groupi_n_1586), .y(csa_tree_add_14_36_groupi_n_1607));
inv csa_tree_add_14_36_groupi_g51342 (.a(csa_tree_add_14_36_groupi_n_1601), .y(csa_tree_add_14_36_groupi_n_1602));
nand2 csa_tree_add_14_36_groupi_g51344__4296 (.a(csa_tree_add_14_36_groupi_n_1561), .b(csa_tree_add_14_36_groupi_n_1501), .y(csa_tree_add_14_36_groupi_n_1599));
nor2 csa_tree_add_14_36_groupi_g51345__3772 (.a(csa_tree_add_14_36_groupi_n_1496), .b(csa_tree_add_14_36_groupi_n_1560), .y(csa_tree_add_14_36_groupi_n_1598));
nand2 csa_tree_add_14_36_groupi_g51346__1474 (.a(csa_tree_add_14_36_groupi_n_1543), .b(csa_tree_add_14_36_groupi_n_1441), .y(csa_tree_add_14_36_groupi_n_1597));
nand2 csa_tree_add_14_36_groupi_g51347__4547 (.a(csa_tree_add_14_36_groupi_n_1474), .b(csa_tree_add_14_36_groupi_n_1552), .y(csa_tree_add_14_36_groupi_n_1596));
nor2 csa_tree_add_14_36_groupi_g51348__9682 (.a(csa_tree_add_14_36_groupi_n_1543), .b(csa_tree_add_14_36_groupi_n_1441), .y(csa_tree_add_14_36_groupi_n_1595));
nand2 csa_tree_add_14_36_groupi_g51349__2683 (.a(csa_tree_add_14_36_groupi_n_1536), .b(csa_tree_add_14_36_groupi_n_2276), .y(csa_tree_add_14_36_groupi_n_1594));
xor2 csa_tree_add_14_36_groupi_g51352__2900 (.a(csa_tree_add_14_36_groupi_n_1484), .b(csa_tree_add_14_36_groupi_n_1356), .y(csa_tree_add_14_36_groupi_n_1591));
nor2 csa_tree_add_14_36_groupi_g51353__2391 (.a(csa_tree_add_14_36_groupi_n_1550), .b(csa_tree_add_14_36_groupi_n_2281), .y(csa_tree_add_14_36_groupi_n_1590));
nand2 csa_tree_add_14_36_groupi_g51354__7675 (.a(csa_tree_add_14_36_groupi_n_1500), .b(csa_tree_add_14_36_groupi_n_2268), .y(csa_tree_add_14_36_groupi_n_1589));
nand2 csa_tree_add_14_36_groupi_g51355__7118 (.a(csa_tree_add_14_36_groupi_n_1540), .b(csa_tree_add_14_36_groupi_n_1512), .y(csa_tree_add_14_36_groupi_n_1588));
nand2 csa_tree_add_14_36_groupi_g51356__8757 (.a(csa_tree_add_14_36_groupi_n_1539), .b(csa_tree_add_14_36_groupi_n_1523), .y(csa_tree_add_14_36_groupi_n_1587));
nand2 csa_tree_add_14_36_groupi_g51357__1786 (.a(csa_tree_add_14_36_groupi_n_2270), .b(csa_tree_add_14_36_groupi_n_2271), .y(csa_tree_add_14_36_groupi_n_1586));
xor2 csa_tree_add_14_36_groupi_g51358__5953 (.a(n_2427), .b(csa_tree_add_14_36_groupi_n_1451), .y(result_0__4_));
xor2 csa_tree_add_14_36_groupi_g51359__5703 (.a(csa_tree_add_14_36_groupi_n_1475), .b(csa_tree_add_14_36_groupi_n_1485), .y(csa_tree_add_14_36_groupi_n_1585));
xor2 csa_tree_add_14_36_groupi_g51360__7114 (.a(csa_tree_add_14_36_groupi_n_1502), .b(csa_tree_add_14_36_groupi_n_1446), .y(csa_tree_add_14_36_groupi_n_1584));
nand2 csa_tree_add_14_36_groupi_g51362__2250 (.a(csa_tree_add_14_36_groupi_n_1316), .b(csa_tree_add_14_36_groupi_n_2130), .y(csa_tree_add_14_36_groupi_n_1605));
xor2 csa_tree_add_14_36_groupi_g51363__6083 (.a(csa_tree_add_14_36_groupi_n_1517), .b(csa_tree_add_14_36_groupi_n_1266), .y(csa_tree_add_14_36_groupi_n_1583));
nand2 csa_tree_add_14_36_groupi_g51364__2703 (.a(csa_tree_add_14_36_groupi_n_2091), .b(csa_tree_add_14_36_groupi_n_1566), .y(csa_tree_add_14_36_groupi_n_1604));
xor2 csa_tree_add_14_36_groupi_g51365__5795 (.a(csa_tree_add_14_36_groupi_n_1497), .b(n_2547), .y(csa_tree_add_14_36_groupi_n_1582));
nor2 csa_tree_add_14_36_groupi_g51366__7344 (.a(csa_tree_add_14_36_groupi_n_2307), .b(csa_tree_add_14_36_groupi_n_1567), .y(csa_tree_add_14_36_groupi_n_1581));
xor2 csa_tree_add_14_36_groupi_g51367__1840 (.a(csa_tree_add_14_36_groupi_n_1494), .b(csa_tree_add_14_36_groupi_n_1441), .y(csa_tree_add_14_36_groupi_n_1580));
nor2 csa_tree_add_14_36_groupi_g51368__5019 (.a(csa_tree_add_14_36_groupi_n_65), .b(csa_tree_add_14_36_groupi_n_2138), .y(csa_tree_add_14_36_groupi_n_1579));
xor2 csa_tree_add_14_36_groupi_g51369__1857 (.a(csa_tree_add_14_36_groupi_n_1492), .b(csa_tree_add_14_36_groupi_n_1471), .y(csa_tree_add_14_36_groupi_n_1578));
nand2 csa_tree_add_14_36_groupi_g51371__8780 (.a(n_2430), .b(n_2429), .y(csa_tree_add_14_36_groupi_n_1601));
xor2 csa_tree_add_14_36_groupi_g51372__4296 (.a(csa_tree_add_14_36_groupi_n_1493), .b(csa_tree_add_14_36_groupi_n_1077), .y(csa_tree_add_14_36_groupi_n_1577));
nand2 csa_tree_add_14_36_groupi_g51374__3772 (.a(csa_tree_add_14_36_groupi_n_1564), .b(csa_tree_add_14_36_groupi_n_2262), .y(csa_tree_add_14_36_groupi_n_1600));
inv csa_tree_add_14_36_groupi_g51376 (.a(csa_tree_add_14_36_groupi_n_1574), .y(csa_tree_add_14_36_groupi_n_1575));
inv csa_tree_add_14_36_groupi_g51377 (.a(csa_tree_add_14_36_groupi_n_2223), .y(csa_tree_add_14_36_groupi_n_1573));
inv csa_tree_add_14_36_groupi_g51378 (.a(csa_tree_add_14_36_groupi_n_1571), .y(csa_tree_add_14_36_groupi_n_1572));
inv csa_tree_add_14_36_groupi_g51380 (.a(csa_tree_add_14_36_groupi_n_2138), .y(csa_tree_add_14_36_groupi_n_1567));
inv csa_tree_add_14_36_groupi_g51381 (.a(csa_tree_add_14_36_groupi_n_2130), .y(csa_tree_add_14_36_groupi_n_1566));
nand2 csa_tree_add_14_36_groupi_g51382__1474 (.a(csa_tree_add_14_36_groupi_n_1525), .b(csa_tree_add_14_36_groupi_n_1468), .y(csa_tree_add_14_36_groupi_n_1565));
nand2 csa_tree_add_14_36_groupi_g51384__4547 (.a(csa_tree_add_14_36_groupi_n_2292), .b(csa_tree_add_14_36_groupi_n_2264), .y(csa_tree_add_14_36_groupi_n_1564));
nand2 csa_tree_add_14_36_groupi_g51385__9682 (.a(csa_tree_add_14_36_groupi_n_1491), .b(csa_tree_add_14_36_groupi_n_1290), .y(csa_tree_add_14_36_groupi_n_1563));
nand2 csa_tree_add_14_36_groupi_g51386__2683 (.a(csa_tree_add_14_36_groupi_n_1504), .b(csa_tree_add_14_36_groupi_n_1466), .y(csa_tree_add_14_36_groupi_n_1562));
nand2 csa_tree_add_14_36_groupi_g51387__1309 (.a(csa_tree_add_14_36_groupi_n_1495), .b(csa_tree_add_14_36_groupi_n_2279), .y(csa_tree_add_14_36_groupi_n_1561));
nor2 csa_tree_add_14_36_groupi_g51388__6877 (.a(csa_tree_add_14_36_groupi_n_1493), .b(csa_tree_add_14_36_groupi_n_1077), .y(csa_tree_add_14_36_groupi_n_1560));
nand2 csa_tree_add_14_36_groupi_g51389__2900 (.a(csa_tree_add_14_36_groupi_n_1493), .b(csa_tree_add_14_36_groupi_n_1077), .y(csa_tree_add_14_36_groupi_n_1559));
nand2 csa_tree_add_14_36_groupi_g51390__2391 (.a(csa_tree_add_14_36_groupi_n_2278), .b(csa_tree_add_14_36_groupi_n_1256), .y(csa_tree_add_14_36_groupi_n_1558));
nand2 csa_tree_add_14_36_groupi_g51391__7675 (.a(csa_tree_add_14_36_groupi_n_1505), .b(csa_tree_add_14_36_groupi_n_1380), .y(csa_tree_add_14_36_groupi_n_1557));
nor2 csa_tree_add_14_36_groupi_g51392__7118 (.a(csa_tree_add_14_36_groupi_n_1514), .b(n_2621), .y(csa_tree_add_14_36_groupi_n_1556));
nor2 csa_tree_add_14_36_groupi_g51393__8757 (.a(csa_tree_add_14_36_groupi_n_2291), .b(csa_tree_add_14_36_groupi_n_1257), .y(csa_tree_add_14_36_groupi_n_1555));
nand2 csa_tree_add_14_36_groupi_g51394__1786 (.a(csa_tree_add_14_36_groupi_n_1489), .b(csa_tree_add_14_36_groupi_n_1406), .y(csa_tree_add_14_36_groupi_n_1554));
nor2 csa_tree_add_14_36_groupi_g51396__5953 (.a(csa_tree_add_14_36_groupi_n_1499), .b(csa_tree_add_14_36_groupi_n_2120), .y(csa_tree_add_14_36_groupi_n_1574));
nor2 csa_tree_add_14_36_groupi_g51398__5703 (.a(csa_tree_add_14_36_groupi_n_1508), .b(csa_tree_add_14_36_groupi_n_1365), .y(csa_tree_add_14_36_groupi_n_1571));
nor2 csa_tree_add_14_36_groupi_g51400__5266 (.a(csa_tree_add_14_36_groupi_n_1381), .b(csa_tree_add_14_36_groupi_n_1509), .y(csa_tree_add_14_36_groupi_n_1569));
nand2 csa_tree_add_14_36_groupi_g51401__2250 (.a(csa_tree_add_14_36_groupi_n_1499), .b(csa_tree_add_14_36_groupi_n_2120), .y(csa_tree_add_14_36_groupi_n_1568));
nand2 csa_tree_add_14_36_groupi_g51403__6083 (.a(csa_tree_add_14_36_groupi_n_1503), .b(csa_tree_add_14_36_groupi_n_1450), .y(csa_tree_add_14_36_groupi_n_2270));
nand2 csa_tree_add_14_36_groupi_g51404__2703 (.a(csa_tree_add_14_36_groupi_n_1517), .b(csa_tree_add_14_36_groupi_n_1267), .y(csa_tree_add_14_36_groupi_n_1553));
nand2 csa_tree_add_14_36_groupi_g51405__5795 (.a(csa_tree_add_14_36_groupi_n_1516), .b(csa_tree_add_14_36_groupi_n_1266), .y(csa_tree_add_14_36_groupi_n_1552));
inv csa_tree_add_14_36_groupi_g51409 (.a(csa_tree_add_14_36_groupi_n_1541), .y(csa_tree_add_14_36_groupi_n_1551));
inv csa_tree_add_14_36_groupi_g51410 (.a(csa_tree_add_14_36_groupi_n_1537), .y(csa_tree_add_14_36_groupi_n_1550));
inv csa_tree_add_14_36_groupi_g51411 (.a(csa_tree_add_14_36_groupi_n_2416), .y(csa_tree_add_14_36_groupi_n_1549));
inv csa_tree_add_14_36_groupi_g51412 (.a(csa_tree_add_14_36_groupi_n_1547), .y(csa_tree_add_14_36_groupi_n_1548));
nor2 csa_tree_add_14_36_groupi_g51414__7344 (.a(csa_tree_add_14_36_groupi_n_1492), .b(csa_tree_add_14_36_groupi_n_1471), .y(csa_tree_add_14_36_groupi_n_1541));
nand2 csa_tree_add_14_36_groupi_g51415__1840 (.a(csa_tree_add_14_36_groupi_n_1492), .b(csa_tree_add_14_36_groupi_n_1471), .y(csa_tree_add_14_36_groupi_n_1540));
xor2 csa_tree_add_14_36_groupi_g51416__5019 (.a(n_2760), .b(csa_tree_add_14_36_groupi_n_1420), .y(result_0__3_));
nand2 csa_tree_add_14_36_groupi_g51417__1857 (.a(csa_tree_add_14_36_groupi_n_1359), .b(csa_tree_add_14_36_groupi_n_1522), .y(csa_tree_add_14_36_groupi_n_1539));
nand2 csa_tree_add_14_36_groupi_g51418__9906 (.a(csa_tree_add_14_36_groupi_n_2277), .b(csa_tree_add_14_36_groupi_n_1255), .y(csa_tree_add_14_36_groupi_n_1538));
nand2 csa_tree_add_14_36_groupi_g51419__8780 (.a(csa_tree_add_14_36_groupi_n_2283), .b(csa_tree_add_14_36_groupi_n_2282), .y(csa_tree_add_14_36_groupi_n_1537));
nand2 csa_tree_add_14_36_groupi_g51420__4296 (.a(csa_tree_add_14_36_groupi_n_1513), .b(csa_tree_add_14_36_groupi_n_2275), .y(csa_tree_add_14_36_groupi_n_1536));
xor2 csa_tree_add_14_36_groupi_g51421__3772 (.a(csa_tree_add_14_36_groupi_n_1186), .b(csa_tree_add_14_36_groupi_n_1428), .y(csa_tree_add_14_36_groupi_n_1535));
xor2 csa_tree_add_14_36_groupi_g51422__1474 (.a(csa_tree_add_14_36_groupi_n_1254), .b(csa_tree_add_14_36_groupi_n_1425), .y(csa_tree_add_14_36_groupi_n_1534));
xor2 csa_tree_add_14_36_groupi_g51423__4547 (.a(csa_tree_add_14_36_groupi_n_1193), .b(csa_tree_add_14_36_groupi_n_1431), .y(csa_tree_add_14_36_groupi_n_1533));
nor2 csa_tree_add_14_36_groupi_g51424__9682 (.a(csa_tree_add_14_36_groupi_n_2283), .b(csa_tree_add_14_36_groupi_n_2282), .y(csa_tree_add_14_36_groupi_n_1532));
xor2 csa_tree_add_14_36_groupi_g51425__2683 (.a(csa_tree_add_14_36_groupi_n_1473), .b(csa_tree_add_14_36_groupi_n_1452), .y(csa_tree_add_14_36_groupi_n_1531));
xor2 csa_tree_add_14_36_groupi_g51426__1309 (.a(csa_tree_add_14_36_groupi_n_1252), .b(csa_tree_add_14_36_groupi_n_1418), .y(csa_tree_add_14_36_groupi_n_1530));
xor2 csa_tree_add_14_36_groupi_g51427__6877 (.a(csa_tree_add_14_36_groupi_n_1476), .b(csa_tree_add_14_36_groupi_n_1432), .y(csa_tree_add_14_36_groupi_n_1529));
xor2 csa_tree_add_14_36_groupi_g51428__2900 (.a(csa_tree_add_14_36_groupi_n_1210), .b(csa_tree_add_14_36_groupi_n_1430), .y(csa_tree_add_14_36_groupi_n_1528));
nand2 csa_tree_add_14_36_groupi_g51429__2391 (.a(csa_tree_add_14_36_groupi_n_1523), .b(csa_tree_add_14_36_groupi_n_1522), .y(csa_tree_add_14_36_groupi_n_1527));
xor2 csa_tree_add_14_36_groupi_g51430__7675 (.a(csa_tree_add_14_36_groupi_n_1429), .b(csa_tree_add_14_36_groupi_n_1214), .y(csa_tree_add_14_36_groupi_n_2416));
xor2 csa_tree_add_14_36_groupi_g51431__7118 (.a(csa_tree_add_14_36_groupi_n_1181), .b(csa_tree_add_14_36_groupi_n_1423), .y(csa_tree_add_14_36_groupi_n_1547));
xor2 csa_tree_add_14_36_groupi_g51433__1786 (.a(csa_tree_add_14_36_groupi_n_1442), .b(csa_tree_add_14_36_groupi_n_1424), .y(csa_tree_add_14_36_groupi_n_2281));
xor2 csa_tree_add_14_36_groupi_g51434__5953 (.a(csa_tree_add_14_36_groupi_n_1247), .b(csa_tree_add_14_36_groupi_n_1421), .y(csa_tree_add_14_36_groupi_n_2268));
xor2 csa_tree_add_14_36_groupi_g51435__5703 (.a(csa_tree_add_14_36_groupi_n_2311), .b(csa_tree_add_14_36_groupi_n_2097), .y(csa_tree_add_14_36_groupi_n_1526));
xor2 csa_tree_add_14_36_groupi_g51438__2250 (.a(csa_tree_add_14_36_groupi_n_1083), .b(csa_tree_add_14_36_groupi_n_1422), .y(csa_tree_add_14_36_groupi_n_2287));
xor2 csa_tree_add_14_36_groupi_g51440__2703 (.a(csa_tree_add_14_36_groupi_n_1355), .b(csa_tree_add_14_36_groupi_n_43), .y(csa_tree_add_14_36_groupi_n_1543));
xor2 csa_tree_add_14_36_groupi_g51441__5795 (.a(csa_tree_add_14_36_groupi_n_1419), .b(n_2561), .y(csa_tree_add_14_36_groupi_n_1542));
inv csa_tree_add_14_36_groupi_g51442 (.a(csa_tree_add_14_36_groupi_n_1506), .y(csa_tree_add_14_36_groupi_n_1525));
inv csa_tree_add_14_36_groupi_g51443 (.a(csa_tree_add_14_36_groupi_n_2176), .y(csa_tree_add_14_36_groupi_n_1524));
inv csa_tree_add_14_36_groupi_g51444 (.a(csa_tree_add_14_36_groupi_n_2255), .y(csa_tree_add_14_36_groupi_n_1521));
inv csa_tree_add_14_36_groupi_g51445 (.a(csa_tree_add_14_36_groupi_n_1519), .y(csa_tree_add_14_36_groupi_n_1520));
inv csa_tree_add_14_36_groupi_g51446 (.a(csa_tree_add_14_36_groupi_n_1517), .y(csa_tree_add_14_36_groupi_n_1516));
inv csa_tree_add_14_36_groupi_g51447 (.a(csa_tree_add_14_36_groupi_n_2291), .y(csa_tree_add_14_36_groupi_n_1514));
inv csa_tree_add_14_36_groupi_g51448 (.a(csa_tree_add_14_36_groupi_n_2277), .y(csa_tree_add_14_36_groupi_n_1513));
nand2 csa_tree_add_14_36_groupi_g51449__7344 (.a(csa_tree_add_14_36_groupi_n_1479), .b(csa_tree_add_14_36_groupi_n_1392), .y(csa_tree_add_14_36_groupi_n_1510));
nor2 csa_tree_add_14_36_groupi_g51450__1840 (.a(csa_tree_add_14_36_groupi_n_1460), .b(csa_tree_add_14_36_groupi_n_1444), .y(csa_tree_add_14_36_groupi_n_1509));
nor2 csa_tree_add_14_36_groupi_g51451__5019 (.a(csa_tree_add_14_36_groupi_n_1442), .b(csa_tree_add_14_36_groupi_n_1368), .y(csa_tree_add_14_36_groupi_n_1508));
nand2 csa_tree_add_14_36_groupi_g51452__1857 (.a(csa_tree_add_14_36_groupi_n_1457), .b(csa_tree_add_14_36_groupi_n_1371), .y(csa_tree_add_14_36_groupi_n_1507));
nor2 csa_tree_add_14_36_groupi_g51454__9906 (.a(csa_tree_add_14_36_groupi_n_1475), .b(csa_tree_add_14_36_groupi_n_1467), .y(csa_tree_add_14_36_groupi_n_1506));
nand2 csa_tree_add_14_36_groupi_g51455__8780 (.a(csa_tree_add_14_36_groupi_n_1473), .b(csa_tree_add_14_36_groupi_n_1379), .y(csa_tree_add_14_36_groupi_n_1505));
nand2 csa_tree_add_14_36_groupi_g51456__4296 (.a(csa_tree_add_14_36_groupi_n_1481), .b(csa_tree_add_14_36_groupi_n_1356), .y(csa_tree_add_14_36_groupi_n_1504));
nand2 csa_tree_add_14_36_groupi_g51457__3772 (.a(csa_tree_add_14_36_groupi_n_1453), .b(csa_tree_add_14_36_groupi_n_1446), .y(csa_tree_add_14_36_groupi_n_1503));
nand2 csa_tree_add_14_36_groupi_g51459__1474 (.a(csa_tree_add_14_36_groupi_n_1447), .b(csa_tree_add_14_36_groupi_n_1315), .y(csa_tree_add_14_36_groupi_n_1523));
nand2 csa_tree_add_14_36_groupi_g51460__4547 (.a(csa_tree_add_14_36_groupi_n_1448), .b(csa_tree_add_14_36_groupi_n_2117), .y(csa_tree_add_14_36_groupi_n_1522));
nor2 csa_tree_add_14_36_groupi_g51462__9682 (.a(csa_tree_add_14_36_groupi_n_1456), .b(csa_tree_add_14_36_groupi_n_1378), .y(csa_tree_add_14_36_groupi_n_1519));
nand2 csa_tree_add_14_36_groupi_g51463__2683 (.a(csa_tree_add_14_36_groupi_n_1458), .b(csa_tree_add_14_36_groupi_n_1397), .y(csa_tree_add_14_36_groupi_n_1518));
nand2 csa_tree_add_14_36_groupi_g51464__1309 (.a(csa_tree_add_14_36_groupi_n_1470), .b(csa_tree_add_14_36_groupi_n_1387), .y(csa_tree_add_14_36_groupi_n_1517));
xor2 csa_tree_add_14_36_groupi_g51465__6877 (.a(csa_tree_add_14_36_groupi_n_1373), .b(csa_tree_add_14_36_groupi_n_582), .y(csa_tree_add_14_36_groupi_n_1502));
nand2 csa_tree_add_14_36_groupi_g51467__2391 (.a(csa_tree_add_14_36_groupi_n_1461), .b(csa_tree_add_14_36_groupi_n_1389), .y(csa_tree_add_14_36_groupi_n_2291));
nand2 csa_tree_add_14_36_groupi_g51468__7675 (.a(csa_tree_add_14_36_groupi_n_1459), .b(csa_tree_add_14_36_groupi_n_1399), .y(csa_tree_add_14_36_groupi_n_2283));
nand2 csa_tree_add_14_36_groupi_g51469__7118 (.a(csa_tree_add_14_36_groupi_n_1464), .b(csa_tree_add_14_36_groupi_n_1386), .y(csa_tree_add_14_36_groupi_n_2277));
nand2 csa_tree_add_14_36_groupi_g51470__8757 (.a(csa_tree_add_14_36_groupi_n_1455), .b(csa_tree_add_14_36_groupi_n_1376), .y(csa_tree_add_14_36_groupi_n_1512));
inv csa_tree_add_14_36_groupi_g51473 (.a(csa_tree_add_14_36_groupi_n_1501), .y(csa_tree_add_14_36_groupi_n_2280));
inv csa_tree_add_14_36_groupi_g51474 (.a(csa_tree_add_14_36_groupi_n_2267), .y(csa_tree_add_14_36_groupi_n_1500));
inv csa_tree_add_14_36_groupi_g51475 (.a(csa_tree_add_14_36_groupi_n_2278), .y(csa_tree_add_14_36_groupi_n_1495));
nand2 csa_tree_add_14_36_groupi_g51476__5953 (.a(csa_tree_add_14_36_groupi_n_1445), .b(csa_tree_add_14_36_groupi_n_1319), .y(csa_tree_add_14_36_groupi_n_1491));
xor2 csa_tree_add_14_36_groupi_g51477__5703 (.a(csa_tree_add_14_36_groupi_n_1339), .b(csa_tree_add_14_36_groupi_n_1076), .y(csa_tree_add_14_36_groupi_n_1490));
nand2 csa_tree_add_14_36_groupi_g51478__7114 (.a(csa_tree_add_14_36_groupi_n_1477), .b(csa_tree_add_14_36_groupi_n_1405), .y(csa_tree_add_14_36_groupi_n_1489));
xor2 csa_tree_add_14_36_groupi_g51479__5266 (.a(csa_tree_add_14_36_groupi_n_1340), .b(n_2768), .y(csa_tree_add_14_36_groupi_n_1488));
nand2 csa_tree_add_14_36_groupi_g51480__2250 (.a(csa_tree_add_14_36_groupi_n_1438), .b(csa_tree_add_14_36_groupi_n_1364), .y(csa_tree_add_14_36_groupi_n_1487));
nand2 csa_tree_add_14_36_groupi_g51481__6083 (.a(csa_tree_add_14_36_groupi_n_1439), .b(csa_tree_add_14_36_groupi_n_1362), .y(csa_tree_add_14_36_groupi_n_1486));
nor2 csa_tree_add_14_36_groupi_g51482__2703 (.a(csa_tree_add_14_36_groupi_n_1434), .b(csa_tree_add_14_36_groupi_n_1383), .y(csa_tree_add_14_36_groupi_n_1501));
nand2 csa_tree_add_14_36_groupi_g51483__5795 (.a(csa_tree_add_14_36_groupi_n_45), .b(csa_tree_add_14_36_groupi_n_1351), .y(csa_tree_add_14_36_groupi_n_2267));
xor2 csa_tree_add_14_36_groupi_g51484__7344 (.a(csa_tree_add_14_36_groupi_n_1185), .b(csa_tree_add_14_36_groupi_n_1330), .y(csa_tree_add_14_36_groupi_n_2292));
xor2 csa_tree_add_14_36_groupi_g51485__1840 (.a(csa_tree_add_14_36_groupi_n_2146), .b(csa_tree_add_14_36_groupi_n_2121), .y(csa_tree_add_14_36_groupi_n_1485));
xor2 csa_tree_add_14_36_groupi_g51486__5019 (.a(n_2609), .b(csa_tree_add_14_36_groupi_n_1227), .y(csa_tree_add_14_36_groupi_n_2271));
xor2 csa_tree_add_14_36_groupi_g51487__1857 (.a(csa_tree_add_14_36_groupi_n_1354), .b(csa_tree_add_14_36_groupi_n_2048), .y(csa_tree_add_14_36_groupi_n_1484));
xor2 csa_tree_add_14_36_groupi_g51488__9906 (.a(csa_tree_add_14_36_groupi_n_1081), .b(csa_tree_add_14_36_groupi_n_1333), .y(csa_tree_add_14_36_groupi_n_1499));
nand2 csa_tree_add_14_36_groupi_g51489__8780 (.a(csa_tree_add_14_36_groupi_n_2311), .b(csa_tree_add_14_36_groupi_n_1478), .y(csa_tree_add_14_36_groupi_n_1483));
nand2 csa_tree_add_14_36_groupi_g51490__4296 (.a(csa_tree_add_14_36_groupi_n_85), .b(csa_tree_add_14_36_groupi_n_2097), .y(csa_tree_add_14_36_groupi_n_1482));
nand2 csa_tree_add_14_36_groupi_g51491__3772 (.a(csa_tree_add_14_36_groupi_n_1437), .b(csa_tree_add_14_36_groupi_n_1374), .y(csa_tree_add_14_36_groupi_n_1498));
xor2 csa_tree_add_14_36_groupi_g51492__1474 (.a(csa_tree_add_14_36_groupi_n_1178), .b(csa_tree_add_14_36_groupi_n_1334), .y(csa_tree_add_14_36_groupi_n_2288));
xor2 csa_tree_add_14_36_groupi_g51493__4547 (.a(csa_tree_add_14_36_groupi_n_1179), .b(csa_tree_add_14_36_groupi_n_1341), .y(csa_tree_add_14_36_groupi_n_2282));
xor2 csa_tree_add_14_36_groupi_g51494__9682 (.a(csa_tree_add_14_36_groupi_n_1085), .b(csa_tree_add_14_36_groupi_n_1332), .y(csa_tree_add_14_36_groupi_n_1497));
nand2 csa_tree_add_14_36_groupi_g51495__2683 (.a(csa_tree_add_14_36_groupi_n_1480), .b(csa_tree_add_14_36_groupi_n_1384), .y(csa_tree_add_14_36_groupi_n_1496));
xor2 csa_tree_add_14_36_groupi_g51496__1309 (.a(csa_tree_add_14_36_groupi_n_1184), .b(csa_tree_add_14_36_groupi_n_1331), .y(csa_tree_add_14_36_groupi_n_2278));
xor2 csa_tree_add_14_36_groupi_g51497__6877 (.a(csa_tree_add_14_36_groupi_n_1191), .b(csa_tree_add_14_36_groupi_n_1337), .y(csa_tree_add_14_36_groupi_n_1494));
xor2 csa_tree_add_14_36_groupi_g51498__2900 (.a(csa_tree_add_14_36_groupi_n_1188), .b(csa_tree_add_14_36_groupi_n_1335), .y(csa_tree_add_14_36_groupi_n_1493));
xor2 csa_tree_add_14_36_groupi_g51499__2391 (.a(csa_tree_add_14_36_groupi_n_1336), .b(n_2556), .y(csa_tree_add_14_36_groupi_n_1492));
inv csa_tree_add_14_36_groupi_g51500 (.a(csa_tree_add_14_36_groupi_n_1465), .y(csa_tree_add_14_36_groupi_n_1481));
inv csa_tree_add_14_36_groupi_g51501 (.a(csa_tree_add_14_36_groupi_n_1463), .y(csa_tree_add_14_36_groupi_n_1480));
inv csa_tree_add_14_36_groupi_g51502 (.a(csa_tree_add_14_36_groupi_n_1462), .y(csa_tree_add_14_36_groupi_n_1479));
inv csa_tree_add_14_36_groupi_g51503 (.a(csa_tree_add_14_36_groupi_n_2097), .y(csa_tree_add_14_36_groupi_n_1478));
inv csa_tree_add_14_36_groupi_g51504 (.a(csa_tree_add_14_36_groupi_n_1476), .y(csa_tree_add_14_36_groupi_n_1477));
nand2 csa_tree_add_14_36_groupi_g51507__7675 (.a(csa_tree_add_14_36_groupi_n_1083), .b(csa_tree_add_14_36_groupi_n_1414), .y(csa_tree_add_14_36_groupi_n_1470));
nand2 csa_tree_add_14_36_groupi_g51509__8757 (.a(csa_tree_add_14_36_groupi_n_2146), .b(csa_tree_add_14_36_groupi_n_2121), .y(csa_tree_add_14_36_groupi_n_1468));
nor2 csa_tree_add_14_36_groupi_g51510__1786 (.a(csa_tree_add_14_36_groupi_n_2146), .b(csa_tree_add_14_36_groupi_n_2121), .y(csa_tree_add_14_36_groupi_n_1467));
nand2 csa_tree_add_14_36_groupi_g51511__5953 (.a(csa_tree_add_14_36_groupi_n_1354), .b(csa_tree_add_14_36_groupi_n_2048), .y(csa_tree_add_14_36_groupi_n_1466));
nor2 csa_tree_add_14_36_groupi_g51512__5703 (.a(csa_tree_add_14_36_groupi_n_1354), .b(csa_tree_add_14_36_groupi_n_2048), .y(csa_tree_add_14_36_groupi_n_1465));
nand2 csa_tree_add_14_36_groupi_g51513__7114 (.a(csa_tree_add_14_36_groupi_n_1193), .b(csa_tree_add_14_36_groupi_n_1412), .y(csa_tree_add_14_36_groupi_n_1464));
nor2 csa_tree_add_14_36_groupi_g51514__5266 (.a(csa_tree_add_14_36_groupi_n_1393), .b(csa_tree_add_14_36_groupi_n_2285), .y(csa_tree_add_14_36_groupi_n_1463));
nor2 csa_tree_add_14_36_groupi_g51515__2250 (.a(csa_tree_add_14_36_groupi_n_2269), .b(csa_tree_add_14_36_groupi_n_1391), .y(csa_tree_add_14_36_groupi_n_1462));
nand2 csa_tree_add_14_36_groupi_g51516__6083 (.a(csa_tree_add_14_36_groupi_n_1415), .b(csa_tree_add_14_36_groupi_n_1132), .y(csa_tree_add_14_36_groupi_n_1461));
nor2 csa_tree_add_14_36_groupi_g51517__2703 (.a(csa_tree_add_14_36_groupi_n_1398), .b(csa_tree_add_14_36_groupi_n_1236), .y(csa_tree_add_14_36_groupi_n_1460));
nand2 csa_tree_add_14_36_groupi_g51518__5795 (.a(csa_tree_add_14_36_groupi_n_1252), .b(csa_tree_add_14_36_groupi_n_1416), .y(csa_tree_add_14_36_groupi_n_1459));
nand2 csa_tree_add_14_36_groupi_g51519__7344 (.a(csa_tree_add_14_36_groupi_n_1417), .b(csa_tree_add_14_36_groupi_n_1177), .y(csa_tree_add_14_36_groupi_n_1458));
nand2 csa_tree_add_14_36_groupi_g51520__1840 (.a(csa_tree_add_14_36_groupi_n_1370), .b(csa_tree_add_14_36_groupi_n_1190), .y(csa_tree_add_14_36_groupi_n_1457));
nor2 csa_tree_add_14_36_groupi_g51521__5019 (.a(csa_tree_add_14_36_groupi_n_1377), .b(csa_tree_add_14_36_groupi_n_1133), .y(csa_tree_add_14_36_groupi_n_1456));
nand2 csa_tree_add_14_36_groupi_g51522__1857 (.a(csa_tree_add_14_36_groupi_n_1211), .b(csa_tree_add_14_36_groupi_n_1375), .y(csa_tree_add_14_36_groupi_n_1455));
nand2 csa_tree_add_14_36_groupi_g51524__8780 (.a(csa_tree_add_14_36_groupi_n_1413), .b(csa_tree_add_14_36_groupi_n_1302), .y(csa_tree_add_14_36_groupi_n_2286));
nand2 csa_tree_add_14_36_groupi_g51526__4296 (.a(csa_tree_add_14_36_groupi_n_1372), .b(csa_tree_add_14_36_groupi_n_582), .y(csa_tree_add_14_36_groupi_n_1453));
xor2 csa_tree_add_14_36_groupi_g51527__3772 (.a(csa_tree_add_14_36_groupi_n_1260), .b(csa_tree_add_14_36_groupi_n_2132), .y(csa_tree_add_14_36_groupi_n_1452));
nand2 csa_tree_add_14_36_groupi_g51528__1474 (.a(csa_tree_add_14_36_groupi_n_1358), .b(csa_tree_add_14_36_groupi_n_1361), .y(csa_tree_add_14_36_groupi_n_1451));
nand2 csa_tree_add_14_36_groupi_g51529__4547 (.a(csa_tree_add_14_36_groupi_n_1373), .b(csa_tree_add_14_36_groupi_n_583), .y(csa_tree_add_14_36_groupi_n_1450));
nand2 csa_tree_add_14_36_groupi_g51530__9682 (.a(csa_tree_add_14_36_groupi_n_1401), .b(csa_tree_add_14_36_groupi_n_1243), .y(csa_tree_add_14_36_groupi_n_1476));
nor2 csa_tree_add_14_36_groupi_g51531__2683 (.a(csa_tree_add_14_36_groupi_n_1347), .b(csa_tree_add_14_36_groupi_n_1281), .y(csa_tree_add_14_36_groupi_n_1475));
nand2 csa_tree_add_14_36_groupi_g51532__1309 (.a(csa_tree_add_14_36_groupi_n_1345), .b(csa_tree_add_14_36_groupi_n_1294), .y(csa_tree_add_14_36_groupi_n_1474));
nand2 csa_tree_add_14_36_groupi_g51533__6877 (.a(csa_tree_add_14_36_groupi_n_1353), .b(csa_tree_add_14_36_groupi_n_1299), .y(csa_tree_add_14_36_groupi_n_1473));
nand2 csa_tree_add_14_36_groupi_g51534__2900 (.a(csa_tree_add_14_36_groupi_n_1402), .b(csa_tree_add_14_36_groupi_n_1301), .y(csa_tree_add_14_36_groupi_n_1472));
nand2 csa_tree_add_14_36_groupi_g51535__2391 (.a(csa_tree_add_14_36_groupi_n_1400), .b(csa_tree_add_14_36_groupi_n_1304), .y(csa_tree_add_14_36_groupi_n_1471));
inv csa_tree_add_14_36_groupi_g51536 (.a(csa_tree_add_14_36_groupi_n_1433), .y(csa_tree_add_14_36_groupi_n_1449));
inv csa_tree_add_14_36_groupi_g51537 (.a(csa_tree_add_14_36_groupi_n_1447), .y(csa_tree_add_14_36_groupi_n_1448));
inv csa_tree_add_14_36_groupi_g51538 (.a(n_2565), .y(csa_tree_add_14_36_groupi_n_1444));
xor2 csa_tree_add_14_36_groupi_g51539__7675 (.a(n_2761), .b(csa_tree_add_14_36_groupi_n_1232), .y(result_0__2_));
xor2 csa_tree_add_14_36_groupi_g51540__7118 (.a(csa_tree_add_14_36_groupi_n_1212), .b(csa_tree_add_14_36_groupi_n_1228), .y(csa_tree_add_14_36_groupi_n_1440));
nand2 csa_tree_add_14_36_groupi_g51541__8757 (.a(csa_tree_add_14_36_groupi_n_1355), .b(csa_tree_add_14_36_groupi_n_1363), .y(csa_tree_add_14_36_groupi_n_1439));
nand2 csa_tree_add_14_36_groupi_g51542__1786 (.a(csa_tree_add_14_36_groupi_n_1187), .b(csa_tree_add_14_36_groupi_n_1369), .y(csa_tree_add_14_36_groupi_n_1438));
nand2 csa_tree_add_14_36_groupi_g51543__5953 (.a(csa_tree_add_14_36_groupi_n_1342), .b(csa_tree_add_14_36_groupi_n_1215), .y(csa_tree_add_14_36_groupi_n_1437));
xor2 csa_tree_add_14_36_groupi_g51545__5703 (.a(csa_tree_add_14_36_groupi_n_1229), .b(n_2614), .y(csa_tree_add_14_36_groupi_n_1436));
xor2 csa_tree_add_14_36_groupi_g51546__7114 (.a(csa_tree_add_14_36_groupi_n_1231), .b(csa_tree_add_14_36_groupi_n_1209), .y(csa_tree_add_14_36_groupi_n_1435));
nor2 csa_tree_add_14_36_groupi_g51547__5266 (.a(csa_tree_add_14_36_groupi_n_1253), .b(csa_tree_add_14_36_groupi_n_1411), .y(csa_tree_add_14_36_groupi_n_1434));
xor2 csa_tree_add_14_36_groupi_g51549__2250 (.a(csa_tree_add_14_36_groupi_n_1259), .b(csa_tree_add_14_36_groupi_n_903), .y(csa_tree_add_14_36_groupi_n_1433));
nand2 csa_tree_add_14_36_groupi_g51550__6083 (.a(csa_tree_add_14_36_groupi_n_1406), .b(csa_tree_add_14_36_groupi_n_1405), .y(csa_tree_add_14_36_groupi_n_1432));
xor2 csa_tree_add_14_36_groupi_g51551__2703 (.a(csa_tree_add_14_36_groupi_n_2101), .b(csa_tree_add_14_36_groupi_n_2067), .y(csa_tree_add_14_36_groupi_n_1431));
xor2 csa_tree_add_14_36_groupi_g51552__5795 (.a(csa_tree_add_14_36_groupi_n_1270), .b(csa_tree_add_14_36_groupi_n_2109), .y(csa_tree_add_14_36_groupi_n_1430));
xor2 csa_tree_add_14_36_groupi_g51553__7344 (.a(csa_tree_add_14_36_groupi_n_1024), .b(csa_tree_add_14_36_groupi_n_1265), .y(csa_tree_add_14_36_groupi_n_1429));
nand2 csa_tree_add_14_36_groupi_g51554__1840 (.a(csa_tree_add_14_36_groupi_n_1364), .b(csa_tree_add_14_36_groupi_n_1369), .y(csa_tree_add_14_36_groupi_n_1428));
xor2 csa_tree_add_14_36_groupi_g51555__5019 (.a(csa_tree_add_14_36_groupi_n_1230), .b(csa_tree_add_14_36_groupi_n_2111), .y(csa_tree_add_14_36_groupi_n_1447));
nand2 csa_tree_add_14_36_groupi_g51556__1857 (.a(csa_tree_add_14_36_groupi_n_1371), .b(csa_tree_add_14_36_groupi_n_1370), .y(csa_tree_add_14_36_groupi_n_1427));
xor2 csa_tree_add_14_36_groupi_g51558__8780 (.a(csa_tree_add_14_36_groupi_n_2151), .b(csa_tree_add_14_36_groupi_n_2095), .y(csa_tree_add_14_36_groupi_n_1425));
nand2 csa_tree_add_14_36_groupi_g51559__4296 (.a(csa_tree_add_14_36_groupi_n_1367), .b(csa_tree_add_14_36_groupi_n_1366), .y(csa_tree_add_14_36_groupi_n_1424));
xor2 csa_tree_add_14_36_groupi_g51560__3772 (.a(csa_tree_add_14_36_groupi_n_1079), .b(csa_tree_add_14_36_groupi_n_1249), .y(csa_tree_add_14_36_groupi_n_1423));
xor2 csa_tree_add_14_36_groupi_g51561__1474 (.a(csa_tree_add_14_36_groupi_n_2093), .b(csa_tree_add_14_36_groupi_n_2037), .y(csa_tree_add_14_36_groupi_n_1422));
xor2 csa_tree_add_14_36_groupi_g51562__4547 (.a(csa_tree_add_14_36_groupi_n_1177), .b(csa_tree_add_14_36_groupi_n_1250), .y(csa_tree_add_14_36_groupi_n_1421));
nand2 csa_tree_add_14_36_groupi_g51563__9682 (.a(csa_tree_add_14_36_groupi_n_1408), .b(n_2425), .y(csa_tree_add_14_36_groupi_n_1420));
xor2 csa_tree_add_14_36_groupi_g51564__2683 (.a(csa_tree_add_14_36_groupi_n_1132), .b(csa_tree_add_14_36_groupi_n_2119), .y(csa_tree_add_14_36_groupi_n_1419));
xor2 csa_tree_add_14_36_groupi_g51565__1309 (.a(csa_tree_add_14_36_groupi_n_1248), .b(csa_tree_add_14_36_groupi_n_2148), .y(csa_tree_add_14_36_groupi_n_1418));
nand2 csa_tree_add_14_36_groupi_g51566__6877 (.a(csa_tree_add_14_36_groupi_n_1349), .b(csa_tree_add_14_36_groupi_n_1286), .y(csa_tree_add_14_36_groupi_n_1446));
nand2 csa_tree_add_14_36_groupi_g51567__2900 (.a(csa_tree_add_14_36_groupi_n_1344), .b(csa_tree_add_14_36_groupi_n_1291), .y(csa_tree_add_14_36_groupi_n_1445));
nand2 csa_tree_add_14_36_groupi_g51569__7675 (.a(csa_tree_add_14_36_groupi_n_1346), .b(csa_tree_add_14_36_groupi_n_1242), .y(csa_tree_add_14_36_groupi_n_1442));
nand2 csa_tree_add_14_36_groupi_g51570__7118 (.a(csa_tree_add_14_36_groupi_n_1343), .b(csa_tree_add_14_36_groupi_n_1287), .y(csa_tree_add_14_36_groupi_n_1441));
inv csa_tree_add_14_36_groupi_g51571 (.a(csa_tree_add_14_36_groupi_n_1396), .y(csa_tree_add_14_36_groupi_n_1417));
inv csa_tree_add_14_36_groupi_g51572 (.a(csa_tree_add_14_36_groupi_n_1395), .y(csa_tree_add_14_36_groupi_n_1416));
inv csa_tree_add_14_36_groupi_g51573 (.a(n_2641), .y(csa_tree_add_14_36_groupi_n_1415));
inv csa_tree_add_14_36_groupi_g51574 (.a(csa_tree_add_14_36_groupi_n_1390), .y(csa_tree_add_14_36_groupi_n_1414));
inv csa_tree_add_14_36_groupi_g51575 (.a(csa_tree_add_14_36_groupi_n_1388), .y(csa_tree_add_14_36_groupi_n_1413));
inv csa_tree_add_14_36_groupi_g51576 (.a(csa_tree_add_14_36_groupi_n_1385), .y(csa_tree_add_14_36_groupi_n_1412));
inv csa_tree_add_14_36_groupi_g51577 (.a(csa_tree_add_14_36_groupi_n_1382), .y(csa_tree_add_14_36_groupi_n_1411));
inv csa_tree_add_14_36_groupi_g51579 (.a(csa_tree_add_14_36_groupi_n_1407), .y(csa_tree_add_14_36_groupi_n_1408));
nand2 csa_tree_add_14_36_groupi_g51581__8757 (.a(csa_tree_add_14_36_groupi_n_1325), .b(n_153), .y(csa_tree_add_14_36_groupi_n_1402));
nand2 csa_tree_add_14_36_groupi_g51583__1786 (.a(csa_tree_add_14_36_groupi_n_1282), .b(csa_tree_add_14_36_groupi_n_1023), .y(csa_tree_add_14_36_groupi_n_1401));
nand2 csa_tree_add_14_36_groupi_g51584__5953 (.a(csa_tree_add_14_36_groupi_n_1081), .b(csa_tree_add_14_36_groupi_n_1326), .y(csa_tree_add_14_36_groupi_n_1400));
nand2 csa_tree_add_14_36_groupi_g51585__5703 (.a(csa_tree_add_14_36_groupi_n_1248), .b(csa_tree_add_14_36_groupi_n_2148), .y(csa_tree_add_14_36_groupi_n_1399));
nand2 csa_tree_add_14_36_groupi_g51586__7114 (.a(csa_tree_add_14_36_groupi_n_1309), .b(csa_tree_add_14_36_groupi_n_1121), .y(csa_tree_add_14_36_groupi_n_1398));
nand2 csa_tree_add_14_36_groupi_g51587__5266 (.a(csa_tree_add_14_36_groupi_n_1247), .b(csa_tree_add_14_36_groupi_n_1250), .y(csa_tree_add_14_36_groupi_n_1397));
nor2 csa_tree_add_14_36_groupi_g51588__2250 (.a(csa_tree_add_14_36_groupi_n_1247), .b(csa_tree_add_14_36_groupi_n_1250), .y(csa_tree_add_14_36_groupi_n_1396));
nor2 csa_tree_add_14_36_groupi_g51589__6083 (.a(csa_tree_add_14_36_groupi_n_1248), .b(csa_tree_add_14_36_groupi_n_2148), .y(csa_tree_add_14_36_groupi_n_1395));
nor2 csa_tree_add_14_36_groupi_g51591__5795 (.a(csa_tree_add_14_36_groupi_n_1192), .b(csa_tree_add_14_36_groupi_n_2300), .y(csa_tree_add_14_36_groupi_n_1393));
nand2 csa_tree_add_14_36_groupi_g51592__7344 (.a(csa_tree_add_14_36_groupi_n_2301), .b(csa_tree_add_14_36_groupi_n_2299), .y(csa_tree_add_14_36_groupi_n_1392));
nor2 csa_tree_add_14_36_groupi_g51593__1840 (.a(csa_tree_add_14_36_groupi_n_2301), .b(csa_tree_add_14_36_groupi_n_2299), .y(csa_tree_add_14_36_groupi_n_1391));
nor2 csa_tree_add_14_36_groupi_g51594__5019 (.a(csa_tree_add_14_36_groupi_n_2093), .b(csa_tree_add_14_36_groupi_n_2037), .y(csa_tree_add_14_36_groupi_n_1390));
nand2 csa_tree_add_14_36_groupi_g51595__1857 (.a(n_2561), .b(csa_tree_add_14_36_groupi_n_2119), .y(csa_tree_add_14_36_groupi_n_1389));
nor2 csa_tree_add_14_36_groupi_g51596__9906 (.a(csa_tree_add_14_36_groupi_n_1191), .b(csa_tree_add_14_36_groupi_n_1296), .y(csa_tree_add_14_36_groupi_n_1388));
nand2 csa_tree_add_14_36_groupi_g51597__8780 (.a(csa_tree_add_14_36_groupi_n_2093), .b(csa_tree_add_14_36_groupi_n_2037), .y(csa_tree_add_14_36_groupi_n_1387));
nand2 csa_tree_add_14_36_groupi_g51598__4296 (.a(csa_tree_add_14_36_groupi_n_2101), .b(csa_tree_add_14_36_groupi_n_2067), .y(csa_tree_add_14_36_groupi_n_1386));
nor2 csa_tree_add_14_36_groupi_g51599__3772 (.a(csa_tree_add_14_36_groupi_n_2101), .b(csa_tree_add_14_36_groupi_n_2067), .y(csa_tree_add_14_36_groupi_n_1385));
nand2 csa_tree_add_14_36_groupi_g51600__1474 (.a(csa_tree_add_14_36_groupi_n_1192), .b(csa_tree_add_14_36_groupi_n_2300), .y(csa_tree_add_14_36_groupi_n_1384));
nor2 csa_tree_add_14_36_groupi_g51601__4547 (.a(csa_tree_add_14_36_groupi_n_2151), .b(csa_tree_add_14_36_groupi_n_2095), .y(csa_tree_add_14_36_groupi_n_1383));
nand2 csa_tree_add_14_36_groupi_g51602__9682 (.a(csa_tree_add_14_36_groupi_n_2151), .b(csa_tree_add_14_36_groupi_n_2095), .y(csa_tree_add_14_36_groupi_n_1382));
nor2 csa_tree_add_14_36_groupi_g51604__2683 (.a(n_2564), .b(csa_tree_add_14_36_groupi_n_1276), .y(csa_tree_add_14_36_groupi_n_1381));
nand2 csa_tree_add_14_36_groupi_g51605__1309 (.a(csa_tree_add_14_36_groupi_n_1261), .b(csa_tree_add_14_36_groupi_n_2132), .y(csa_tree_add_14_36_groupi_n_1380));
nand2 csa_tree_add_14_36_groupi_g51606__6877 (.a(csa_tree_add_14_36_groupi_n_1260), .b(csa_tree_add_14_36_groupi_n_1142), .y(csa_tree_add_14_36_groupi_n_1379));
nor2 csa_tree_add_14_36_groupi_g51607__2900 (.a(csa_tree_add_14_36_groupi_n_1259), .b(csa_tree_add_14_36_groupi_n_903), .y(csa_tree_add_14_36_groupi_n_1378));
nor2 csa_tree_add_14_36_groupi_g51608__2391 (.a(csa_tree_add_14_36_groupi_n_1258), .b(csa_tree_add_14_36_groupi_n_2061), .y(csa_tree_add_14_36_groupi_n_1377));
nand2 csa_tree_add_14_36_groupi_g51609__7675 (.a(csa_tree_add_14_36_groupi_n_1270), .b(csa_tree_add_14_36_groupi_n_1312), .y(csa_tree_add_14_36_groupi_n_1376));
nand2 csa_tree_add_14_36_groupi_g51610__7118 (.a(csa_tree_add_14_36_groupi_n_1269), .b(csa_tree_add_14_36_groupi_n_2109), .y(csa_tree_add_14_36_groupi_n_1375));
nor2 csa_tree_add_14_36_groupi_g51612__1786 (.a(csa_tree_add_14_36_groupi_n_965), .b(csa_tree_add_14_36_groupi_n_1263), .y(csa_tree_add_14_36_groupi_n_1407));
nand2 csa_tree_add_14_36_groupi_g51613__5953 (.a(csa_tree_add_14_36_groupi_n_1272), .b(csa_tree_add_14_36_groupi_n_1311), .y(csa_tree_add_14_36_groupi_n_1406));
nand2 csa_tree_add_14_36_groupi_g51614__5703 (.a(csa_tree_add_14_36_groupi_n_1273), .b(csa_tree_add_14_36_groupi_n_2104), .y(csa_tree_add_14_36_groupi_n_1405));
nand2 csa_tree_add_14_36_groupi_g51615__7114 (.a(csa_tree_add_14_36_groupi_n_1025), .b(csa_tree_add_14_36_groupi_n_1265), .y(csa_tree_add_14_36_groupi_n_1374));
nand2 csa_tree_add_14_36_groupi_g51618__6083 (.a(csa_tree_add_14_36_groupi_n_1234), .b(csa_tree_add_14_36_groupi_n_1197), .y(csa_tree_add_14_36_groupi_n_1403));
inv csa_tree_add_14_36_groupi_g51622 (.a(csa_tree_add_14_36_groupi_n_1372), .y(csa_tree_add_14_36_groupi_n_1373));
inv csa_tree_add_14_36_groupi_g51623 (.a(csa_tree_add_14_36_groupi_n_1367), .y(csa_tree_add_14_36_groupi_n_1368));
inv csa_tree_add_14_36_groupi_g51624 (.a(csa_tree_add_14_36_groupi_n_1365), .y(csa_tree_add_14_36_groupi_n_1366));
inv csa_tree_add_14_36_groupi_g51627 (.a(n_2434), .y(csa_tree_add_14_36_groupi_n_1361));
inv csa_tree_add_14_36_groupi_g51628 (.a(csa_tree_add_14_36_groupi_n_1358), .y(csa_tree_add_14_36_groupi_n_1357));
nand2 csa_tree_add_14_36_groupi_g51629__2703 (.a(csa_tree_add_14_36_groupi_n_1184), .b(csa_tree_add_14_36_groupi_n_1321), .y(csa_tree_add_14_36_groupi_n_1353));
nor2 csa_tree_add_14_36_groupi_g51630__5795 (.a(csa_tree_add_14_36_groupi_n_1079), .b(csa_tree_add_14_36_groupi_n_1249), .y(csa_tree_add_14_36_groupi_n_1352));
nand2 csa_tree_add_14_36_groupi_g51631__7344 (.a(csa_tree_add_14_36_groupi_n_1079), .b(csa_tree_add_14_36_groupi_n_1249), .y(csa_tree_add_14_36_groupi_n_1351));
nand2 csa_tree_add_14_36_groupi_g51632__1840 (.a(csa_tree_add_14_36_groupi_n_1283), .b(csa_tree_add_14_36_groupi_n_1139), .y(csa_tree_add_14_36_groupi_n_1350));
nand2 csa_tree_add_14_36_groupi_g51633__5019 (.a(csa_tree_add_14_36_groupi_n_1188), .b(csa_tree_add_14_36_groupi_n_1329), .y(csa_tree_add_14_36_groupi_n_1349));
nor2 csa_tree_add_14_36_groupi_g51635__9906 (.a(csa_tree_add_14_36_groupi_n_1180), .b(csa_tree_add_14_36_groupi_n_1278), .y(csa_tree_add_14_36_groupi_n_1347));
nand2 csa_tree_add_14_36_groupi_g51636__8780 (.a(csa_tree_add_14_36_groupi_n_1284), .b(csa_tree_add_14_36_groupi_n_1137), .y(csa_tree_add_14_36_groupi_n_1346));
nand2 csa_tree_add_14_36_groupi_g51637__4296 (.a(csa_tree_add_14_36_groupi_n_1178), .b(csa_tree_add_14_36_groupi_n_1320), .y(csa_tree_add_14_36_groupi_n_1345));
nand2 csa_tree_add_14_36_groupi_g51638__3772 (.a(csa_tree_add_14_36_groupi_n_1185), .b(csa_tree_add_14_36_groupi_n_1327), .y(csa_tree_add_14_36_groupi_n_1344));
nand2 csa_tree_add_14_36_groupi_g51639__1474 (.a(csa_tree_add_14_36_groupi_n_1085), .b(csa_tree_add_14_36_groupi_n_1322), .y(csa_tree_add_14_36_groupi_n_1343));
xor2 csa_tree_add_14_36_groupi_g51640__4547 (.a(n_2642), .b(csa_tree_add_14_36_groupi_n_1065), .y(csa_tree_add_14_36_groupi_n_1372));
nand2 csa_tree_add_14_36_groupi_g51641__9682 (.a(csa_tree_add_14_36_groupi_n_1274), .b(csa_tree_add_14_36_groupi_n_1222), .y(csa_tree_add_14_36_groupi_n_1371));
nand2 csa_tree_add_14_36_groupi_g51642__2683 (.a(csa_tree_add_14_36_groupi_n_1275), .b(csa_tree_add_14_36_groupi_n_2122), .y(csa_tree_add_14_36_groupi_n_1370));
nand2 csa_tree_add_14_36_groupi_g51643__1309 (.a(csa_tree_add_14_36_groupi_n_1090), .b(csa_tree_add_14_36_groupi_n_2152), .y(csa_tree_add_14_36_groupi_n_2264));
nand2 csa_tree_add_14_36_groupi_g51644__6877 (.a(csa_tree_add_14_36_groupi_n_1089), .b(csa_tree_add_14_36_groupi_n_1318), .y(csa_tree_add_14_36_groupi_n_2262));
nand2 csa_tree_add_14_36_groupi_g51645__2900 (.a(csa_tree_add_14_36_groupi_n_2114), .b(csa_tree_add_14_36_groupi_n_1313), .y(csa_tree_add_14_36_groupi_n_1369));
nand2 csa_tree_add_14_36_groupi_g51646__2391 (.a(csa_tree_add_14_36_groupi_n_1262), .b(csa_tree_add_14_36_groupi_n_2118), .y(csa_tree_add_14_36_groupi_n_1367));
nor2 csa_tree_add_14_36_groupi_g51647__7675 (.a(csa_tree_add_14_36_groupi_n_1262), .b(csa_tree_add_14_36_groupi_n_2118), .y(csa_tree_add_14_36_groupi_n_1365));
nand2 csa_tree_add_14_36_groupi_g51648__7118 (.a(csa_tree_add_14_36_groupi_n_1219), .b(csa_tree_add_14_36_groupi_n_2113), .y(csa_tree_add_14_36_groupi_n_1364));
nand2 csa_tree_add_14_36_groupi_g51649__8757 (.a(csa_tree_add_14_36_groupi_n_1024), .b(csa_tree_add_14_36_groupi_n_1264), .y(csa_tree_add_14_36_groupi_n_1342));
nand2 csa_tree_add_14_36_groupi_g51650__1786 (.a(csa_tree_add_14_36_groupi_n_2088), .b(csa_tree_add_14_36_groupi_n_1317), .y(csa_tree_add_14_36_groupi_n_1363));
nand2 csa_tree_add_14_36_groupi_g51651__5953 (.a(csa_tree_add_14_36_groupi_n_1314), .b(csa_tree_add_14_36_groupi_n_2099), .y(csa_tree_add_14_36_groupi_n_1362));
nand2 csa_tree_add_14_36_groupi_g51652__5703 (.a(csa_tree_add_14_36_groupi_n_1280), .b(csa_tree_add_14_36_groupi_n_1279), .y(csa_tree_add_14_36_groupi_n_1341));
xor2 csa_tree_add_14_36_groupi_g51653__7114 (.a(n_2765), .b(n_2762), .y(csa_tree_add_14_36_groupi_n_1340));
xor2 csa_tree_add_14_36_groupi_g51654__5266 (.a(csa_tree_add_14_36_groupi_n_1139), .b(csa_tree_add_14_36_groupi_n_1175), .y(csa_tree_add_14_36_groupi_n_1339));
xor2 csa_tree_add_14_36_groupi_g51656__6083 (.a(csa_tree_add_14_36_groupi_n_1174), .b(csa_tree_add_14_36_groupi_n_1078), .y(csa_tree_add_14_36_groupi_n_1338));
xor2 csa_tree_add_14_36_groupi_g51657__2703 (.a(csa_tree_add_14_36_groupi_n_1075), .b(csa_tree_add_14_36_groupi_n_2046), .y(csa_tree_add_14_36_groupi_n_1337));
xor2 csa_tree_add_14_36_groupi_g51658__5795 (.a(csa_tree_add_14_36_groupi_n_1023), .b(csa_tree_add_14_36_groupi_n_2108), .y(csa_tree_add_14_36_groupi_n_1336));
xor2 csa_tree_add_14_36_groupi_g51659__7344 (.a(csa_tree_add_14_36_groupi_n_2096), .b(csa_tree_add_14_36_groupi_n_2107), .y(csa_tree_add_14_36_groupi_n_1335));
xor2 csa_tree_add_14_36_groupi_g51660__1840 (.a(csa_tree_add_14_36_groupi_n_2125), .b(csa_tree_add_14_36_groupi_n_2133), .y(csa_tree_add_14_36_groupi_n_1334));
xor2 csa_tree_add_14_36_groupi_g51661__5019 (.a(csa_tree_add_14_36_groupi_n_2058), .b(csa_tree_add_14_36_groupi_n_2147), .y(csa_tree_add_14_36_groupi_n_1333));
xor2 csa_tree_add_14_36_groupi_g51662__1857 (.a(csa_tree_add_14_36_groupi_n_2090), .b(csa_tree_add_14_36_groupi_n_2126), .y(csa_tree_add_14_36_groupi_n_1332));
xor2 csa_tree_add_14_36_groupi_g51663__9906 (.a(csa_tree_add_14_36_groupi_n_2150), .b(csa_tree_add_14_36_groupi_n_2100), .y(csa_tree_add_14_36_groupi_n_1331));
xor2 csa_tree_add_14_36_groupi_g51664__8780 (.a(csa_tree_add_14_36_groupi_n_2042), .b(csa_tree_add_14_36_groupi_n_2112), .y(csa_tree_add_14_36_groupi_n_1330));
nand2 csa_tree_add_14_36_groupi_g51665__4296 (.a(csa_tree_add_14_36_groupi_n_1237), .b(csa_tree_add_14_36_groupi_n_1198), .y(csa_tree_add_14_36_groupi_n_1359));
nand2 csa_tree_add_14_36_groupi_g51666__3772 (.a(n_2432), .b(n_2433), .y(csa_tree_add_14_36_groupi_n_1358));
nand2 csa_tree_add_14_36_groupi_g51667__1474 (.a(csa_tree_add_14_36_groupi_n_1245), .b(csa_tree_add_14_36_groupi_n_1202), .y(csa_tree_add_14_36_groupi_n_1356));
nand2 csa_tree_add_14_36_groupi_g51668__4547 (.a(n_2778), .b(csa_tree_add_14_36_groupi_n_1002), .y(csa_tree_add_14_36_groupi_n_1355));
xor2 csa_tree_add_14_36_groupi_g51669__9682 (.a(n_2781), .b(csa_tree_add_14_36_groupi_n_1054), .y(csa_tree_add_14_36_groupi_n_1354));
inv csa_tree_add_14_36_groupi_g51670 (.a(csa_tree_add_14_36_groupi_n_1308), .y(csa_tree_add_14_36_groupi_n_1329));
inv csa_tree_add_14_36_groupi_g51672 (.a(csa_tree_add_14_36_groupi_n_1305), .y(csa_tree_add_14_36_groupi_n_1327));
inv csa_tree_add_14_36_groupi_g51673 (.a(csa_tree_add_14_36_groupi_n_1303), .y(csa_tree_add_14_36_groupi_n_1326));
inv csa_tree_add_14_36_groupi_g51674 (.a(csa_tree_add_14_36_groupi_n_1300), .y(csa_tree_add_14_36_groupi_n_1325));
inv csa_tree_add_14_36_groupi_g51677 (.a(csa_tree_add_14_36_groupi_n_1295), .y(csa_tree_add_14_36_groupi_n_1322));
inv csa_tree_add_14_36_groupi_g51678 (.a(csa_tree_add_14_36_groupi_n_1293), .y(csa_tree_add_14_36_groupi_n_1321));
inv csa_tree_add_14_36_groupi_g51679 (.a(csa_tree_add_14_36_groupi_n_1292), .y(csa_tree_add_14_36_groupi_n_1320));
inv csa_tree_add_14_36_groupi_g51680 (.a(csa_tree_add_14_36_groupi_n_1289), .y(csa_tree_add_14_36_groupi_n_1319));
inv csa_tree_add_14_36_groupi_g51681 (.a(csa_tree_add_14_36_groupi_n_2152), .y(csa_tree_add_14_36_groupi_n_1318));
inv csa_tree_add_14_36_groupi_g51682 (.a(csa_tree_add_14_36_groupi_n_2099), .y(csa_tree_add_14_36_groupi_n_1317));
inv csa_tree_add_14_36_groupi_g51683 (.a(csa_tree_add_14_36_groupi_n_2091), .y(csa_tree_add_14_36_groupi_n_1316));
inv csa_tree_add_14_36_groupi_g51684 (.a(csa_tree_add_14_36_groupi_n_2117), .y(csa_tree_add_14_36_groupi_n_1315));
inv csa_tree_add_14_36_groupi_g51685 (.a(csa_tree_add_14_36_groupi_n_2088), .y(csa_tree_add_14_36_groupi_n_1314));
inv csa_tree_add_14_36_groupi_g51686 (.a(csa_tree_add_14_36_groupi_n_2113), .y(csa_tree_add_14_36_groupi_n_1313));
inv csa_tree_add_14_36_groupi_g51687 (.a(csa_tree_add_14_36_groupi_n_2109), .y(csa_tree_add_14_36_groupi_n_1312));
inv csa_tree_add_14_36_groupi_g51688 (.a(csa_tree_add_14_36_groupi_n_2104), .y(csa_tree_add_14_36_groupi_n_1311));
nor2 csa_tree_add_14_36_groupi_g51689__2683 (.a(csa_tree_add_14_36_groupi_n_1217), .b(csa_tree_add_14_36_groupi_n_1029), .y(csa_tree_add_14_36_groupi_n_1309));
nor2 csa_tree_add_14_36_groupi_g51690__1309 (.a(csa_tree_add_14_36_groupi_n_2096), .b(csa_tree_add_14_36_groupi_n_2107), .y(csa_tree_add_14_36_groupi_n_1308));
nor2 csa_tree_add_14_36_groupi_g51693__2391 (.a(csa_tree_add_14_36_groupi_n_2042), .b(csa_tree_add_14_36_groupi_n_2112), .y(csa_tree_add_14_36_groupi_n_1305));
nand2 csa_tree_add_14_36_groupi_g51694__7675 (.a(csa_tree_add_14_36_groupi_n_2058), .b(csa_tree_add_14_36_groupi_n_2147), .y(csa_tree_add_14_36_groupi_n_1304));
nor2 csa_tree_add_14_36_groupi_g51695__7118 (.a(csa_tree_add_14_36_groupi_n_2058), .b(csa_tree_add_14_36_groupi_n_2147), .y(csa_tree_add_14_36_groupi_n_1303));
nand2 csa_tree_add_14_36_groupi_g51696__8757 (.a(csa_tree_add_14_36_groupi_n_1075), .b(csa_tree_add_14_36_groupi_n_2046), .y(csa_tree_add_14_36_groupi_n_1302));
nand2 csa_tree_add_14_36_groupi_g51697__1786 (.a(csa_tree_add_14_36_groupi_n_2131), .b(csa_tree_add_14_36_groupi_n_2111), .y(csa_tree_add_14_36_groupi_n_1301));
nor2 csa_tree_add_14_36_groupi_g51698__5953 (.a(csa_tree_add_14_36_groupi_n_2131), .b(csa_tree_add_14_36_groupi_n_2111), .y(csa_tree_add_14_36_groupi_n_1300));
nand2 csa_tree_add_14_36_groupi_g51699__5703 (.a(csa_tree_add_14_36_groupi_n_2150), .b(csa_tree_add_14_36_groupi_n_2100), .y(csa_tree_add_14_36_groupi_n_1299));
nor2 csa_tree_add_14_36_groupi_g51702__2250 (.a(csa_tree_add_14_36_groupi_n_1075), .b(csa_tree_add_14_36_groupi_n_2046), .y(csa_tree_add_14_36_groupi_n_1296));
nor2 csa_tree_add_14_36_groupi_g51703__6083 (.a(csa_tree_add_14_36_groupi_n_2090), .b(csa_tree_add_14_36_groupi_n_2126), .y(csa_tree_add_14_36_groupi_n_1295));
nand2 csa_tree_add_14_36_groupi_g51704__2703 (.a(csa_tree_add_14_36_groupi_n_2125), .b(csa_tree_add_14_36_groupi_n_2133), .y(csa_tree_add_14_36_groupi_n_1294));
nor2 csa_tree_add_14_36_groupi_g51705__5795 (.a(csa_tree_add_14_36_groupi_n_2150), .b(csa_tree_add_14_36_groupi_n_2100), .y(csa_tree_add_14_36_groupi_n_1293));
nor2 csa_tree_add_14_36_groupi_g51706__7344 (.a(csa_tree_add_14_36_groupi_n_2125), .b(csa_tree_add_14_36_groupi_n_2133), .y(csa_tree_add_14_36_groupi_n_1292));
nand2 csa_tree_add_14_36_groupi_g51707__1840 (.a(csa_tree_add_14_36_groupi_n_2042), .b(csa_tree_add_14_36_groupi_n_2112), .y(csa_tree_add_14_36_groupi_n_1291));
nand2 csa_tree_add_14_36_groupi_g51708__5019 (.a(csa_tree_add_14_36_groupi_n_1174), .b(csa_tree_add_14_36_groupi_n_1078), .y(csa_tree_add_14_36_groupi_n_1290));
nor2 csa_tree_add_14_36_groupi_g51709__1857 (.a(csa_tree_add_14_36_groupi_n_1174), .b(csa_tree_add_14_36_groupi_n_1078), .y(csa_tree_add_14_36_groupi_n_1289));
nand2 csa_tree_add_14_36_groupi_g51710__9906 (.a(csa_tree_add_14_36_groupi_n_1200), .b(csa_tree_add_14_36_groupi_n_1155), .y(csa_tree_add_14_36_groupi_n_1288));
nand2 csa_tree_add_14_36_groupi_g51711__8780 (.a(csa_tree_add_14_36_groupi_n_2090), .b(csa_tree_add_14_36_groupi_n_2126), .y(csa_tree_add_14_36_groupi_n_1287));
nand2 csa_tree_add_14_36_groupi_g51712__4296 (.a(csa_tree_add_14_36_groupi_n_2096), .b(csa_tree_add_14_36_groupi_n_2107), .y(csa_tree_add_14_36_groupi_n_1286));
xor2 csa_tree_add_14_36_groupi_g51717__3772 (.a(csa_tree_add_14_36_groupi_n_1093), .b(csa_tree_add_14_36_groupi_n_2077), .y(csa_tree_add_14_36_groupi_n_1285));
inv csa_tree_add_14_36_groupi_g51734 (.a(n_2658), .y(csa_tree_add_14_36_groupi_n_1284));
inv csa_tree_add_14_36_groupi_g51735 (.a(csa_tree_add_14_36_groupi_n_1238), .y(csa_tree_add_14_36_groupi_n_1283));
inv csa_tree_add_14_36_groupi_g51736 (.a(n_2635), .y(csa_tree_add_14_36_groupi_n_1282));
inv csa_tree_add_14_36_groupi_g51737 (.a(csa_tree_add_14_36_groupi_n_1280), .y(csa_tree_add_14_36_groupi_n_1281));
inv csa_tree_add_14_36_groupi_g51738 (.a(csa_tree_add_14_36_groupi_n_1278), .y(csa_tree_add_14_36_groupi_n_1279));
inv csa_tree_add_14_36_groupi_g51740 (.a(csa_tree_add_14_36_groupi_n_1274), .y(csa_tree_add_14_36_groupi_n_1275));
inv csa_tree_add_14_36_groupi_g51741 (.a(csa_tree_add_14_36_groupi_n_1272), .y(csa_tree_add_14_36_groupi_n_1273));
inv csa_tree_add_14_36_groupi_g51743 (.a(csa_tree_add_14_36_groupi_n_1270), .y(csa_tree_add_14_36_groupi_n_1269));
inv csa_tree_add_14_36_groupi_g51744 (.a(csa_tree_add_14_36_groupi_n_1266), .y(csa_tree_add_14_36_groupi_n_1267));
inv csa_tree_add_14_36_groupi_g51745 (.a(csa_tree_add_14_36_groupi_n_1265), .y(csa_tree_add_14_36_groupi_n_1264));
inv csa_tree_add_14_36_groupi_g51746 (.a(csa_tree_add_14_36_groupi_n_1260), .y(csa_tree_add_14_36_groupi_n_1261));
inv csa_tree_add_14_36_groupi_g51747 (.a(csa_tree_add_14_36_groupi_n_1259), .y(csa_tree_add_14_36_groupi_n_1258));
inv csa_tree_add_14_36_groupi_g51748 (.a(n_2621), .y(csa_tree_add_14_36_groupi_n_1257));
inv csa_tree_add_14_36_groupi_g51749 (.a(csa_tree_add_14_36_groupi_n_2279), .y(csa_tree_add_14_36_groupi_n_1256));
inv csa_tree_add_14_36_groupi_g51750 (.a(csa_tree_add_14_36_groupi_n_2275), .y(csa_tree_add_14_36_groupi_n_1255));
inv csa_tree_add_14_36_groupi_g51751 (.a(csa_tree_add_14_36_groupi_n_1253), .y(csa_tree_add_14_36_groupi_n_1254));
xor2 csa_tree_add_14_36_groupi_g51752__4547 (.a(csa_tree_add_14_36_groupi_n_1138), .b(csa_tree_add_14_36_groupi_n_921), .y(csa_tree_add_14_36_groupi_n_1246));
nand2 csa_tree_add_14_36_groupi_g51753__9682 (.a(csa_tree_add_14_36_groupi_n_1212), .b(csa_tree_add_14_36_groupi_n_1226), .y(csa_tree_add_14_36_groupi_n_1245));
nand2 csa_tree_add_14_36_groupi_g51755__1309 (.a(n_2556), .b(csa_tree_add_14_36_groupi_n_2108), .y(csa_tree_add_14_36_groupi_n_1243));
nand2 csa_tree_add_14_36_groupi_g51756__6877 (.a(n_2614), .b(csa_tree_add_14_36_groupi_n_2128), .y(csa_tree_add_14_36_groupi_n_1242));
nand2 csa_tree_add_14_36_groupi_g51757__2900 (.a(csa_tree_add_14_36_groupi_n_1225), .b(csa_tree_add_14_36_groupi_n_836), .y(csa_tree_add_14_36_groupi_n_1241));
nand2 csa_tree_add_14_36_groupi_g51759__7675 (.a(csa_tree_add_14_36_groupi_n_1076), .b(csa_tree_add_14_36_groupi_n_1175), .y(csa_tree_add_14_36_groupi_n_1239));
nor2 csa_tree_add_14_36_groupi_g51760__7118 (.a(csa_tree_add_14_36_groupi_n_1076), .b(csa_tree_add_14_36_groupi_n_1175), .y(csa_tree_add_14_36_groupi_n_1238));
nand2 csa_tree_add_14_36_groupi_g51761__8757 (.a(csa_tree_add_14_36_groupi_n_1195), .b(csa_tree_add_14_36_groupi_n_1209), .y(csa_tree_add_14_36_groupi_n_1237));
nand2 csa_tree_add_14_36_groupi_g51762__1786 (.a(csa_tree_add_14_36_groupi_n_1154), .b(csa_tree_add_14_36_groupi_n_1223), .y(csa_tree_add_14_36_groupi_n_1236));
xor2 csa_tree_add_14_36_groupi_g51763__5953 (.a(csa_tree_add_14_36_groupi_n_1135), .b(csa_tree_add_14_36_groupi_n_923), .y(csa_tree_add_14_36_groupi_n_1235));
nand2 csa_tree_add_14_36_groupi_g51764__5703 (.a(csa_tree_add_14_36_groupi_n_1196), .b(csa_tree_add_14_36_groupi_n_1216), .y(csa_tree_add_14_36_groupi_n_1234));
nand2 csa_tree_add_14_36_groupi_g51766__5266 (.a(csa_tree_add_14_36_groupi_n_1160), .b(csa_tree_add_14_36_groupi_n_1027), .y(csa_tree_add_14_36_groupi_n_2276));
nor2 csa_tree_add_14_36_groupi_g51767__2250 (.a(csa_tree_add_14_36_groupi_n_1221), .b(n_2759), .y(csa_tree_add_14_36_groupi_n_1232));
nand2 csa_tree_add_14_36_groupi_g51768__6083 (.a(csa_tree_add_14_36_groupi_n_1092), .b(csa_tree_add_14_36_groupi_n_2145), .y(csa_tree_add_14_36_groupi_n_1280));
nor2 csa_tree_add_14_36_groupi_g51769__2703 (.a(csa_tree_add_14_36_groupi_n_1092), .b(csa_tree_add_14_36_groupi_n_2145), .y(csa_tree_add_14_36_groupi_n_1278));
xor2 csa_tree_add_14_36_groupi_g51770__5795 (.a(csa_tree_add_14_36_groupi_n_1141), .b(n_153), .y(csa_tree_add_14_36_groupi_n_1231));
nor2 csa_tree_add_14_36_groupi_g51771__7344 (.a(csa_tree_add_14_36_groupi_n_1217), .b(csa_tree_add_14_36_groupi_n_1224), .y(csa_tree_add_14_36_groupi_n_1276));
xor2 csa_tree_add_14_36_groupi_g51772__1840 (.a(n_2654), .b(csa_tree_add_14_36_groupi_n_1056), .y(csa_tree_add_14_36_groupi_n_1274));
xor2 csa_tree_add_14_36_groupi_g51773__5019 (.a(csa_tree_add_14_36_groupi_n_788), .b(csa_tree_add_14_36_groupi_n_1053), .y(csa_tree_add_14_36_groupi_n_1272));
xor2 csa_tree_add_14_36_groupi_g51775__9906 (.a(n_153), .b(csa_tree_add_14_36_groupi_n_2131), .y(csa_tree_add_14_36_groupi_n_1230));
xor2 csa_tree_add_14_36_groupi_g51776__8780 (.a(n_2631), .b(csa_tree_add_14_36_groupi_n_1049), .y(csa_tree_add_14_36_groupi_n_1270));
xor2 csa_tree_add_14_36_groupi_g51777__4296 (.a(csa_tree_add_14_36_groupi_n_1137), .b(csa_tree_add_14_36_groupi_n_2128), .y(csa_tree_add_14_36_groupi_n_1229));
xor2 csa_tree_add_14_36_groupi_g51779__1474 (.a(csa_tree_add_14_36_groupi_n_1086), .b(csa_tree_add_14_36_groupi_n_1063), .y(csa_tree_add_14_36_groupi_n_1266));
xor2 csa_tree_add_14_36_groupi_g51780__4547 (.a(csa_tree_add_14_36_groupi_n_1080), .b(csa_tree_add_14_36_groupi_n_2105), .y(csa_tree_add_14_36_groupi_n_1228));
xor2 csa_tree_add_14_36_groupi_g51781__9682 (.a(csa_tree_add_14_36_groupi_n_871), .b(csa_tree_add_14_36_groupi_n_1055), .y(csa_tree_add_14_36_groupi_n_1265));
xor2 csa_tree_add_14_36_groupi_g51782__2683 (.a(csa_tree_add_14_36_groupi_n_963), .b(csa_tree_add_14_36_groupi_n_1046), .y(csa_tree_add_14_36_groupi_n_1263));
xor2 csa_tree_add_14_36_groupi_g51783__1309 (.a(csa_tree_add_14_36_groupi_n_1066), .b(csa_tree_add_14_36_groupi_n_2144), .y(csa_tree_add_14_36_groupi_n_2269));
xor2 csa_tree_add_14_36_groupi_g51784__6877 (.a(csa_tree_add_14_36_groupi_n_776), .b(csa_tree_add_14_36_groupi_n_1060), .y(csa_tree_add_14_36_groupi_n_1262));
nand2 csa_tree_add_14_36_groupi_g51785__2900 (.a(csa_tree_add_14_36_groupi_n_1205), .b(csa_tree_add_14_36_groupi_n_1043), .y(csa_tree_add_14_36_groupi_n_1260));
xor2 csa_tree_add_14_36_groupi_g51786__2391 (.a(csa_tree_add_14_36_groupi_n_2272), .b(n_2605), .y(csa_tree_add_14_36_groupi_n_1227));
xor2 csa_tree_add_14_36_groupi_g51787__7675 (.a(csa_tree_add_14_36_groupi_n_872), .b(csa_tree_add_14_36_groupi_n_1051), .y(csa_tree_add_14_36_groupi_n_1259));
xor2 csa_tree_add_14_36_groupi_g51789__8757 (.a(csa_tree_add_14_36_groupi_n_1084), .b(csa_tree_add_14_36_groupi_n_1059), .y(csa_tree_add_14_36_groupi_n_2279));
xor2 csa_tree_add_14_36_groupi_g51790__1786 (.a(csa_tree_add_14_36_groupi_n_1064), .b(csa_tree_add_14_36_groupi_n_2031), .y(csa_tree_add_14_36_groupi_n_2275));
xor2 csa_tree_add_14_36_groupi_g51791__5953 (.a(csa_tree_add_14_36_groupi_n_869), .b(csa_tree_add_14_36_groupi_n_1057), .y(csa_tree_add_14_36_groupi_n_1253));
nand2 csa_tree_add_14_36_groupi_g51792__5703 (.a(csa_tree_add_14_36_groupi_n_1206), .b(csa_tree_add_14_36_groupi_n_1045), .y(csa_tree_add_14_36_groupi_n_1252));
xor2 csa_tree_add_14_36_groupi_g51793__7114 (.a(csa_tree_add_14_36_groupi_n_870), .b(csa_tree_add_14_36_groupi_n_1052), .y(csa_tree_add_14_36_groupi_n_1251));
xor2 csa_tree_add_14_36_groupi_g51794__5266 (.a(csa_tree_add_14_36_groupi_n_964), .b(csa_tree_add_14_36_groupi_n_1062), .y(csa_tree_add_14_36_groupi_n_1250));
xor2 csa_tree_add_14_36_groupi_g51795__2250 (.a(csa_tree_add_14_36_groupi_n_779), .b(csa_tree_add_14_36_groupi_n_1050), .y(csa_tree_add_14_36_groupi_n_1249));
xor2 csa_tree_add_14_36_groupi_g51796__6083 (.a(csa_tree_add_14_36_groupi_n_873), .b(csa_tree_add_14_36_groupi_n_1047), .y(csa_tree_add_14_36_groupi_n_1248));
xor2 csa_tree_add_14_36_groupi_g51797__2703 (.a(csa_tree_add_14_36_groupi_n_1136), .b(csa_tree_add_14_36_groupi_n_1061), .y(csa_tree_add_14_36_groupi_n_1247));
inv csa_tree_add_14_36_groupi_g51798 (.a(csa_tree_add_14_36_groupi_n_1201), .y(csa_tree_add_14_36_groupi_n_1226));
inv csa_tree_add_14_36_groupi_g51799 (.a(csa_tree_add_14_36_groupi_n_1199), .y(csa_tree_add_14_36_groupi_n_1225));
inv csa_tree_add_14_36_groupi_g51800 (.a(csa_tree_add_14_36_groupi_n_1223), .y(csa_tree_add_14_36_groupi_n_1224));
inv csa_tree_add_14_36_groupi_g51801 (.a(csa_tree_add_14_36_groupi_n_2122), .y(csa_tree_add_14_36_groupi_n_1222));
inv csa_tree_add_14_36_groupi_g51802 (.a(n_2753), .y(csa_tree_add_14_36_groupi_n_1221));
inv csa_tree_add_14_36_groupi_g51803 (.a(csa_tree_add_14_36_groupi_n_2114), .y(csa_tree_add_14_36_groupi_n_1219));
inv csa_tree_add_14_36_groupi_g51804 (.a(csa_tree_add_14_36_groupi_n_1214), .y(csa_tree_add_14_36_groupi_n_1215));
inv csa_tree_add_14_36_groupi_g51805 (.a(csa_tree_add_14_36_groupi_n_1210), .y(csa_tree_add_14_36_groupi_n_1211));
nand2 csa_tree_add_14_36_groupi_g51806__5795 (.a(csa_tree_add_14_36_groupi_n_1082), .b(csa_tree_add_14_36_groupi_n_1009), .y(csa_tree_add_14_36_groupi_n_1206));
nand2 csa_tree_add_14_36_groupi_g51807__7344 (.a(csa_tree_add_14_36_groupi_n_1084), .b(csa_tree_add_14_36_groupi_n_1006), .y(csa_tree_add_14_36_groupi_n_1205));
nand2 csa_tree_add_14_36_groupi_g51808__1840 (.a(csa_tree_add_14_36_groupi_n_1087), .b(csa_tree_add_14_36_groupi_n_1038), .y(csa_tree_add_14_36_groupi_n_1204));
nand2 csa_tree_add_14_36_groupi_g51809__5019 (.a(csa_tree_add_14_36_groupi_n_1136), .b(csa_tree_add_14_36_groupi_n_1030), .y(csa_tree_add_14_36_groupi_n_1203));
nand2 csa_tree_add_14_36_groupi_g51810__1857 (.a(csa_tree_add_14_36_groupi_n_1080), .b(csa_tree_add_14_36_groupi_n_2105), .y(csa_tree_add_14_36_groupi_n_1202));
nor2 csa_tree_add_14_36_groupi_g51811__9906 (.a(csa_tree_add_14_36_groupi_n_1080), .b(csa_tree_add_14_36_groupi_n_2105), .y(csa_tree_add_14_36_groupi_n_1201));
nand2 csa_tree_add_14_36_groupi_g51812__8780 (.a(csa_tree_add_14_36_groupi_n_1138), .b(csa_tree_add_14_36_groupi_n_709), .y(csa_tree_add_14_36_groupi_n_1200));
nor2 csa_tree_add_14_36_groupi_g51813__4296 (.a(csa_tree_add_14_36_groupi_n_1135), .b(csa_tree_add_14_36_groupi_n_833), .y(csa_tree_add_14_36_groupi_n_1199));
nand2 csa_tree_add_14_36_groupi_g51814__3772 (.a(csa_tree_add_14_36_groupi_n_1141), .b(csa_tree_add_14_36_groupi_n_81), .y(csa_tree_add_14_36_groupi_n_1198));
nand2 csa_tree_add_14_36_groupi_g51815__1474 (.a(n_2637), .b(csa_tree_add_14_36_groupi_n_1088), .y(csa_tree_add_14_36_groupi_n_1223));
nand2 csa_tree_add_14_36_groupi_g51817__4547 (.a(csa_tree_add_14_36_groupi_n_1094), .b(csa_tree_add_14_36_groupi_n_2077), .y(csa_tree_add_14_36_groupi_n_1197));
nand2 csa_tree_add_14_36_groupi_g51820__2683 (.a(csa_tree_add_14_36_groupi_n_1093), .b(csa_tree_add_14_36_groupi_n_807), .y(csa_tree_add_14_36_groupi_n_1196));
nor2 csa_tree_add_14_36_groupi_g51823__6877 (.a(n_2637), .b(csa_tree_add_14_36_groupi_n_1088), .y(csa_tree_add_14_36_groupi_n_1217));
nand2 csa_tree_add_14_36_groupi_g51824__2900 (.a(csa_tree_add_14_36_groupi_n_1140), .b(n_153), .y(csa_tree_add_14_36_groupi_n_1195));
nand2 csa_tree_add_14_36_groupi_g51825__2391 (.a(csa_tree_add_14_36_groupi_n_1120), .b(csa_tree_add_14_36_groupi_n_1016), .y(csa_tree_add_14_36_groupi_n_1216));
nand2 csa_tree_add_14_36_groupi_g51826__7675 (.a(csa_tree_add_14_36_groupi_n_1118), .b(csa_tree_add_14_36_groupi_n_1015), .y(csa_tree_add_14_36_groupi_n_1214));
nand2 csa_tree_add_14_36_groupi_g51828__8757 (.a(csa_tree_add_14_36_groupi_n_1115), .b(csa_tree_add_14_36_groupi_n_930), .y(csa_tree_add_14_36_groupi_n_1212));
nand2 csa_tree_add_14_36_groupi_g51829__1786 (.a(csa_tree_add_14_36_groupi_n_1149), .b(csa_tree_add_14_36_groupi_n_1012), .y(csa_tree_add_14_36_groupi_n_1210));
nand2 csa_tree_add_14_36_groupi_g51831__5953 (.a(csa_tree_add_14_36_groupi_n_1147), .b(csa_tree_add_14_36_groupi_n_998), .y(csa_tree_add_14_36_groupi_n_1209));
inv csa_tree_add_14_36_groupi_g51847 (.a(csa_tree_add_14_36_groupi_n_1192), .y(csa_tree_add_14_36_groupi_n_2284));
inv csa_tree_add_14_36_groupi_g51848 (.a(csa_tree_add_14_36_groupi_n_1189), .y(csa_tree_add_14_36_groupi_n_1190));
inv csa_tree_add_14_36_groupi_g51849 (.a(csa_tree_add_14_36_groupi_n_1186), .y(csa_tree_add_14_36_groupi_n_1187));
inv csa_tree_add_14_36_groupi_g51851 (.a(csa_tree_add_14_36_groupi_n_1179), .y(csa_tree_add_14_36_groupi_n_1180));
xor2 csa_tree_add_14_36_groupi_g51852__5266 (.a(csa_tree_add_14_36_groupi_n_907), .b(csa_tree_add_14_36_groupi_n_801), .y(csa_tree_add_14_36_groupi_n_1172));
xor2 csa_tree_add_14_36_groupi_g51853__2250 (.a(csa_tree_add_14_36_groupi_n_909), .b(csa_tree_add_14_36_groupi_n_790), .y(csa_tree_add_14_36_groupi_n_1171));
xor2 csa_tree_add_14_36_groupi_g51854__6083 (.a(csa_tree_add_14_36_groupi_n_910), .b(csa_tree_add_14_36_groupi_n_785), .y(csa_tree_add_14_36_groupi_n_1170));
xor2 csa_tree_add_14_36_groupi_g51855__2703 (.a(csa_tree_add_14_36_groupi_n_917), .b(csa_tree_add_14_36_groupi_n_713), .y(csa_tree_add_14_36_groupi_n_1169));
xor2 csa_tree_add_14_36_groupi_g51856__5795 (.a(csa_tree_add_14_36_groupi_n_911), .b(csa_tree_add_14_36_groupi_n_803), .y(csa_tree_add_14_36_groupi_n_1168));
xor2 csa_tree_add_14_36_groupi_g51857__7344 (.a(csa_tree_add_14_36_groupi_n_916), .b(csa_tree_add_14_36_groupi_n_723), .y(csa_tree_add_14_36_groupi_n_1167));
xor2 csa_tree_add_14_36_groupi_g51858__1840 (.a(csa_tree_add_14_36_groupi_n_920), .b(csa_tree_add_14_36_groupi_n_731), .y(csa_tree_add_14_36_groupi_n_1166));
xor2 csa_tree_add_14_36_groupi_g51859__5019 (.a(csa_tree_add_14_36_groupi_n_922), .b(csa_tree_add_14_36_groupi_n_778), .y(csa_tree_add_14_36_groupi_n_1165));
xor2 csa_tree_add_14_36_groupi_g51860__1857 (.a(csa_tree_add_14_36_groupi_n_912), .b(csa_tree_add_14_36_groupi_n_726), .y(csa_tree_add_14_36_groupi_n_1164));
xor2 csa_tree_add_14_36_groupi_g51861__9906 (.a(csa_tree_add_14_36_groupi_n_919), .b(csa_tree_add_14_36_groupi_n_722), .y(csa_tree_add_14_36_groupi_n_1163));
xor2 csa_tree_add_14_36_groupi_g51862__8780 (.a(csa_tree_add_14_36_groupi_n_906), .b(csa_tree_add_14_36_groupi_n_730), .y(csa_tree_add_14_36_groupi_n_1162));
nand2 csa_tree_add_14_36_groupi_g51864__3772 (.a(csa_tree_add_14_36_groupi_n_1086), .b(csa_tree_add_14_36_groupi_n_1031), .y(csa_tree_add_14_36_groupi_n_1160));
nand2 csa_tree_add_14_36_groupi_g51869__1309 (.a(csa_tree_add_14_36_groupi_n_1069), .b(csa_tree_add_14_36_groupi_n_736), .y(csa_tree_add_14_36_groupi_n_1155));
nand2 csa_tree_add_14_36_groupi_g51870__6877 (.a(csa_tree_add_14_36_groupi_n_1122), .b(csa_tree_add_14_36_groupi_n_793), .y(csa_tree_add_14_36_groupi_n_1154));
xor2 csa_tree_add_14_36_groupi_g51871__2900 (.a(csa_tree_add_14_36_groupi_n_905), .b(csa_tree_add_14_36_groupi_n_498), .y(result_0__1_));
xor2 csa_tree_add_14_36_groupi_g51872__2391 (.a(csa_tree_add_14_36_groupi_n_868), .b(csa_tree_add_14_36_groupi_n_908), .y(csa_tree_add_14_36_groupi_n_1153));
xor2 csa_tree_add_14_36_groupi_g51873__7675 (.a(csa_tree_add_14_36_groupi_n_918), .b(csa_tree_add_14_36_groupi_n_727), .y(csa_tree_add_14_36_groupi_n_1152));
xor2 csa_tree_add_14_36_groupi_g51874__7118 (.a(csa_tree_add_14_36_groupi_n_931), .b(csa_tree_add_14_36_groupi_n_729), .y(csa_tree_add_14_36_groupi_n_1151));
nand2 csa_tree_add_14_36_groupi_g51876__1786 (.a(csa_tree_add_14_36_groupi_n_1073), .b(csa_tree_add_14_36_groupi_n_957), .y(csa_tree_add_14_36_groupi_n_1193));
nor2 csa_tree_add_14_36_groupi_g51877__5953 (.a(csa_tree_add_14_36_groupi_n_1072), .b(csa_tree_add_14_36_groupi_n_960), .y(csa_tree_add_14_36_groupi_n_1192));
nor2 csa_tree_add_14_36_groupi_g51878__5703 (.a(csa_tree_add_14_36_groupi_n_1070), .b(csa_tree_add_14_36_groupi_n_969), .y(csa_tree_add_14_36_groupi_n_1191));
nand2 csa_tree_add_14_36_groupi_g51879__7114 (.a(csa_tree_add_14_36_groupi_n_1109), .b(csa_tree_add_14_36_groupi_n_1020), .y(csa_tree_add_14_36_groupi_n_1189));
nand2 csa_tree_add_14_36_groupi_g51880__5266 (.a(csa_tree_add_14_36_groupi_n_1101), .b(csa_tree_add_14_36_groupi_n_974), .y(csa_tree_add_14_36_groupi_n_1188));
nand2 csa_tree_add_14_36_groupi_g51881__2250 (.a(csa_tree_add_14_36_groupi_n_1102), .b(csa_tree_add_14_36_groupi_n_976), .y(csa_tree_add_14_36_groupi_n_1186));
nand2 csa_tree_add_14_36_groupi_g51882__6083 (.a(csa_tree_add_14_36_groupi_n_1106), .b(csa_tree_add_14_36_groupi_n_1026), .y(csa_tree_add_14_36_groupi_n_1185));
nand2 csa_tree_add_14_36_groupi_g51883__2703 (.a(csa_tree_add_14_36_groupi_n_1130), .b(csa_tree_add_14_36_groupi_n_986), .y(csa_tree_add_14_36_groupi_n_1184));
nand2 csa_tree_add_14_36_groupi_g51886__1840 (.a(csa_tree_add_14_36_groupi_n_1148), .b(csa_tree_add_14_36_groupi_n_981), .y(csa_tree_add_14_36_groupi_n_1181));
nand2 csa_tree_add_14_36_groupi_g51887__5019 (.a(csa_tree_add_14_36_groupi_n_1146), .b(csa_tree_add_14_36_groupi_n_994), .y(csa_tree_add_14_36_groupi_n_1179));
nand2 csa_tree_add_14_36_groupi_g51888__1857 (.a(csa_tree_add_14_36_groupi_n_1111), .b(csa_tree_add_14_36_groupi_n_997), .y(csa_tree_add_14_36_groupi_n_1178));
nand2 csa_tree_add_14_36_groupi_g51889__9906 (.a(csa_tree_add_14_36_groupi_n_1144), .b(csa_tree_add_14_36_groupi_n_1018), .y(csa_tree_add_14_36_groupi_n_1177));
xor2 csa_tree_add_14_36_groupi_g51891__4296 (.a(csa_tree_add_14_36_groupi_n_913), .b(csa_tree_add_14_36_groupi_n_721), .y(csa_tree_add_14_36_groupi_n_1175));
nand2 csa_tree_add_14_36_groupi_g51892__3772 (.a(csa_tree_add_14_36_groupi_n_1113), .b(csa_tree_add_14_36_groupi_n_1007), .y(csa_tree_add_14_36_groupi_n_1174));
inv csa_tree_add_14_36_groupi_g51895 (.a(csa_tree_add_14_36_groupi_n_1128), .y(csa_tree_add_14_36_groupi_n_1149));
inv csa_tree_add_14_36_groupi_g51896 (.a(csa_tree_add_14_36_groupi_n_1127), .y(csa_tree_add_14_36_groupi_n_1148));
inv csa_tree_add_14_36_groupi_g51897 (.a(csa_tree_add_14_36_groupi_n_1126), .y(csa_tree_add_14_36_groupi_n_1147));
inv csa_tree_add_14_36_groupi_g51898 (.a(csa_tree_add_14_36_groupi_n_1125), .y(csa_tree_add_14_36_groupi_n_1146));
inv csa_tree_add_14_36_groupi_g51900 (.a(csa_tree_add_14_36_groupi_n_1112), .y(csa_tree_add_14_36_groupi_n_1144));
inv csa_tree_add_14_36_groupi_g51902 (.a(csa_tree_add_14_36_groupi_n_2132), .y(csa_tree_add_14_36_groupi_n_1142));
inv csa_tree_add_14_36_groupi_g51903 (.a(csa_tree_add_14_36_groupi_n_1141), .y(csa_tree_add_14_36_groupi_n_1140));
nand2 csa_tree_add_14_36_groupi_g51904__4547 (.a(csa_tree_add_14_36_groupi_n_869), .b(csa_tree_add_14_36_groupi_n_1034), .y(csa_tree_add_14_36_groupi_n_1130));
nor2 csa_tree_add_14_36_groupi_g51906__2683 (.a(csa_tree_add_14_36_groupi_n_871), .b(csa_tree_add_14_36_groupi_n_983), .y(csa_tree_add_14_36_groupi_n_1128));
nor2 csa_tree_add_14_36_groupi_g51907__1309 (.a(csa_tree_add_14_36_groupi_n_872), .b(csa_tree_add_14_36_groupi_n_992), .y(csa_tree_add_14_36_groupi_n_1127));
nor2 csa_tree_add_14_36_groupi_g51908__6877 (.a(csa_tree_add_14_36_groupi_n_788), .b(csa_tree_add_14_36_groupi_n_999), .y(csa_tree_add_14_36_groupi_n_1126));
nor2 csa_tree_add_14_36_groupi_g51909__2900 (.a(csa_tree_add_14_36_groupi_n_873), .b(csa_tree_add_14_36_groupi_n_993), .y(csa_tree_add_14_36_groupi_n_1125));
nand2 csa_tree_add_14_36_groupi_g51911__7675 (.a(csa_tree_add_14_36_groupi_n_937), .b(csa_tree_add_14_36_groupi_n_820), .y(csa_tree_add_14_36_groupi_n_1123));
nor2 csa_tree_add_14_36_groupi_g51912__7118 (.a(csa_tree_add_14_36_groupi_n_1021), .b(csa_tree_add_14_36_groupi_n_2055), .y(csa_tree_add_14_36_groupi_n_1122));
nand2 csa_tree_add_14_36_groupi_g51913__8757 (.a(csa_tree_add_14_36_groupi_n_800), .b(csa_tree_add_14_36_groupi_n_1022), .y(csa_tree_add_14_36_groupi_n_1121));
nand2 csa_tree_add_14_36_groupi_g51914__1786 (.a(csa_tree_add_14_36_groupi_n_1042), .b(csa_tree_add_14_36_groupi_n_964), .y(csa_tree_add_14_36_groupi_n_1120));
nand2 csa_tree_add_14_36_groupi_g51915__5953 (.a(csa_tree_add_14_36_groupi_n_938), .b(csa_tree_add_14_36_groupi_n_831), .y(csa_tree_add_14_36_groupi_n_1119));
nand2 csa_tree_add_14_36_groupi_g51916__5703 (.a(csa_tree_add_14_36_groupi_n_776), .b(csa_tree_add_14_36_groupi_n_1037), .y(csa_tree_add_14_36_groupi_n_1118));
nand2 csa_tree_add_14_36_groupi_g51918__5266 (.a(csa_tree_add_14_36_groupi_n_941), .b(csa_tree_add_14_36_groupi_n_838), .y(csa_tree_add_14_36_groupi_n_1116));
nand2 csa_tree_add_14_36_groupi_g51919__2250 (.a(csa_tree_add_14_36_groupi_n_924), .b(csa_tree_add_14_36_groupi_n_2144), .y(csa_tree_add_14_36_groupi_n_1115));
nand2 csa_tree_add_14_36_groupi_g51920__6083 (.a(csa_tree_add_14_36_groupi_n_942), .b(csa_tree_add_14_36_groupi_n_842), .y(csa_tree_add_14_36_groupi_n_1114));
nand2 csa_tree_add_14_36_groupi_g51921__2703 (.a(csa_tree_add_14_36_groupi_n_1044), .b(n_147), .y(csa_tree_add_14_36_groupi_n_1113));
nor2 csa_tree_add_14_36_groupi_g51922__5795 (.a(csa_tree_add_14_36_groupi_n_779), .b(csa_tree_add_14_36_groupi_n_984), .y(csa_tree_add_14_36_groupi_n_1112));
nand2 csa_tree_add_14_36_groupi_g51923__7344 (.a(csa_tree_add_14_36_groupi_n_1039), .b(n_127), .y(csa_tree_add_14_36_groupi_n_1111));
nand2 csa_tree_add_14_36_groupi_g51924__1840 (.a(csa_tree_add_14_36_groupi_n_943), .b(csa_tree_add_14_36_groupi_n_843), .y(csa_tree_add_14_36_groupi_n_1110));
nand2 csa_tree_add_14_36_groupi_g51925__5019 (.a(csa_tree_add_14_36_groupi_n_1036), .b(csa_tree_add_14_36_groupi_n_870), .y(csa_tree_add_14_36_groupi_n_1109));
nand2 csa_tree_add_14_36_groupi_g51926__1857 (.a(csa_tree_add_14_36_groupi_n_939), .b(csa_tree_add_14_36_groupi_n_840), .y(csa_tree_add_14_36_groupi_n_1108));
nand2 csa_tree_add_14_36_groupi_g51927__9906 (.a(csa_tree_add_14_36_groupi_n_945), .b(csa_tree_add_14_36_groupi_n_847), .y(csa_tree_add_14_36_groupi_n_1107));
nand2 csa_tree_add_14_36_groupi_g51928__8780 (.a(csa_tree_add_14_36_groupi_n_966), .b(csa_tree_add_14_36_groupi_n_2031), .y(csa_tree_add_14_36_groupi_n_1106));
nand2 csa_tree_add_14_36_groupi_g51929__4296 (.a(csa_tree_add_14_36_groupi_n_946), .b(csa_tree_add_14_36_groupi_n_849), .y(csa_tree_add_14_36_groupi_n_1105));
nand2 csa_tree_add_14_36_groupi_g51930__3772 (.a(csa_tree_add_14_36_groupi_n_1040), .b(csa_tree_add_14_36_groupi_n_963), .y(csa_tree_add_14_36_groupi_n_1104));
nand2 csa_tree_add_14_36_groupi_g51932__4547 (.a(csa_tree_add_14_36_groupi_n_1041), .b(n_149), .y(csa_tree_add_14_36_groupi_n_1102));
nand2 csa_tree_add_14_36_groupi_g51933__9682 (.a(csa_tree_add_14_36_groupi_n_1032), .b(n_139), .y(csa_tree_add_14_36_groupi_n_1101));
nand2 csa_tree_add_14_36_groupi_g51934__2683 (.a(csa_tree_add_14_36_groupi_n_954), .b(csa_tree_add_14_36_groupi_n_845), .y(csa_tree_add_14_36_groupi_n_1100));
nand2 csa_tree_add_14_36_groupi_g51935__1309 (.a(csa_tree_add_14_36_groupi_n_953), .b(csa_tree_add_14_36_groupi_n_865), .y(csa_tree_add_14_36_groupi_n_1099));
nand2 csa_tree_add_14_36_groupi_g51936__6877 (.a(csa_tree_add_14_36_groupi_n_950), .b(csa_tree_add_14_36_groupi_n_857), .y(csa_tree_add_14_36_groupi_n_1098));
nand2 csa_tree_add_14_36_groupi_g51937__2900 (.a(csa_tree_add_14_36_groupi_n_949), .b(csa_tree_add_14_36_groupi_n_859), .y(csa_tree_add_14_36_groupi_n_1097));
nand2 csa_tree_add_14_36_groupi_g51938__2391 (.a(csa_tree_add_14_36_groupi_n_967), .b(csa_tree_add_14_36_groupi_n_855), .y(csa_tree_add_14_36_groupi_n_1096));
nand2 csa_tree_add_14_36_groupi_g51939__7675 (.a(csa_tree_add_14_36_groupi_n_947), .b(csa_tree_add_14_36_groupi_n_851), .y(csa_tree_add_14_36_groupi_n_1095));
nand2 csa_tree_add_14_36_groupi_g51941__7118 (.a(csa_tree_add_14_36_groupi_n_968), .b(csa_tree_add_14_36_groupi_n_412), .y(csa_tree_add_14_36_groupi_n_1141));
nand2 csa_tree_add_14_36_groupi_g51942__8757 (.a(csa_tree_add_14_36_groupi_n_944), .b(csa_tree_add_14_36_groupi_n_844), .y(csa_tree_add_14_36_groupi_n_1139));
nand2 csa_tree_add_14_36_groupi_g51943__1786 (.a(csa_tree_add_14_36_groupi_n_1028), .b(csa_tree_add_14_36_groupi_n_874), .y(csa_tree_add_14_36_groupi_n_1138));
nand2 csa_tree_add_14_36_groupi_g51944__5953 (.a(csa_tree_add_14_36_groupi_n_959), .b(csa_tree_add_14_36_groupi_n_752), .y(csa_tree_add_14_36_groupi_n_1137));
nand2 csa_tree_add_14_36_groupi_g51945__5703 (.a(csa_tree_add_14_36_groupi_n_961), .b(csa_tree_add_14_36_groupi_n_793), .y(csa_tree_add_14_36_groupi_n_1136));
nor2 csa_tree_add_14_36_groupi_g51946__7114 (.a(csa_tree_add_14_36_groupi_n_952), .b(csa_tree_add_14_36_groupi_n_825), .y(csa_tree_add_14_36_groupi_n_1135));
nand2 csa_tree_add_14_36_groupi_g51948__2250 (.a(csa_tree_add_14_36_groupi_n_962), .b(csa_tree_add_14_36_groupi_n_751), .y(csa_tree_add_14_36_groupi_n_1133));
nand2 csa_tree_add_14_36_groupi_g51949__6083 (.a(csa_tree_add_14_36_groupi_n_972), .b(csa_tree_add_14_36_groupi_n_813), .y(csa_tree_add_14_36_groupi_n_1132));
inv csa_tree_add_14_36_groupi_g51952 (.a(csa_tree_add_14_36_groupi_n_1093), .y(csa_tree_add_14_36_groupi_n_1094));
inv csa_tree_add_14_36_groupi_g51953 (.a(csa_tree_add_14_36_groupi_n_1089), .y(csa_tree_add_14_36_groupi_n_1090));
nand2 csa_tree_add_14_36_groupi_g51954__5795 (.a(csa_tree_add_14_36_groupi_n_936), .b(csa_tree_add_14_36_groupi_n_824), .y(csa_tree_add_14_36_groupi_n_1074));
nand2 csa_tree_add_14_36_groupi_g51955__7344 (.a(csa_tree_add_14_36_groupi_n_1017), .b(csa_tree_add_14_36_groupi_n_61), .y(csa_tree_add_14_36_groupi_n_1073));
nor2 csa_tree_add_14_36_groupi_g51956__1840 (.a(csa_tree_add_14_36_groupi_n_970), .b(n_139), .y(csa_tree_add_14_36_groupi_n_1072));
nor2 csa_tree_add_14_36_groupi_g51957__5019 (.a(csa_tree_add_14_36_groupi_n_955), .b(n_145), .y(csa_tree_add_14_36_groupi_n_1071));
nor2 csa_tree_add_14_36_groupi_g51958__1857 (.a(csa_tree_add_14_36_groupi_n_1010), .b(n_127), .y(csa_tree_add_14_36_groupi_n_1070));
nand2 csa_tree_add_14_36_groupi_g51959__9906 (.a(csa_tree_add_14_36_groupi_n_1028), .b(csa_tree_add_14_36_groupi_n_940), .y(csa_tree_add_14_36_groupi_n_1069));
nand2 csa_tree_add_14_36_groupi_g51960__8780 (.a(csa_tree_add_14_36_groupi_n_934), .b(csa_tree_add_14_36_groupi_n_828), .y(csa_tree_add_14_36_groupi_n_1068));
nand2 csa_tree_add_14_36_groupi_g51961__4296 (.a(csa_tree_add_14_36_groupi_n_933), .b(csa_tree_add_14_36_groupi_n_821), .y(csa_tree_add_14_36_groupi_n_1067));
xor2 csa_tree_add_14_36_groupi_g51962__3772 (.a(n_125), .b(csa_tree_add_14_36_groupi_n_2044), .y(csa_tree_add_14_36_groupi_n_1066));
xor2 csa_tree_add_14_36_groupi_g51963__1474 (.a(csa_tree_add_14_36_groupi_n_2140), .b(csa_tree_add_14_36_groupi_n_2092), .y(csa_tree_add_14_36_groupi_n_1065));
nand2 csa_tree_add_14_36_groupi_g51964__4547 (.a(csa_tree_add_14_36_groupi_n_1026), .b(csa_tree_add_14_36_groupi_n_966), .y(csa_tree_add_14_36_groupi_n_1064));
nand2 csa_tree_add_14_36_groupi_g51965__9682 (.a(csa_tree_add_14_36_groupi_n_1027), .b(csa_tree_add_14_36_groupi_n_1031), .y(csa_tree_add_14_36_groupi_n_1063));
xor2 csa_tree_add_14_36_groupi_g51966__2683 (.a(csa_tree_add_14_36_groupi_n_816), .b(csa_tree_add_14_36_groupi_n_2056), .y(csa_tree_add_14_36_groupi_n_1093));
xor2 csa_tree_add_14_36_groupi_g51967__1309 (.a(csa_tree_add_14_36_groupi_n_2072), .b(csa_tree_add_14_36_groupi_n_2050), .y(csa_tree_add_14_36_groupi_n_1062));
xor2 csa_tree_add_14_36_groupi_g51968__6877 (.a(csa_tree_add_14_36_groupi_n_2029), .b(csa_tree_add_14_36_groupi_n_2053), .y(csa_tree_add_14_36_groupi_n_1061));
xor2 csa_tree_add_14_36_groupi_g51969__2900 (.a(csa_tree_add_14_36_groupi_n_2070), .b(csa_tree_add_14_36_groupi_n_2052), .y(csa_tree_add_14_36_groupi_n_1060));
xor2 csa_tree_add_14_36_groupi_g51970__2391 (.a(csa_tree_add_14_36_groupi_n_2038), .b(csa_tree_add_14_36_groupi_n_2045), .y(csa_tree_add_14_36_groupi_n_1059));
xor2 csa_tree_add_14_36_groupi_g51971__7675 (.a(csa_tree_add_14_36_groupi_n_814), .b(csa_tree_add_14_36_groupi_n_2079), .y(csa_tree_add_14_36_groupi_n_1092));
xor2 csa_tree_add_14_36_groupi_g51973__8757 (.a(csa_tree_add_14_36_groupi_n_2083), .b(csa_tree_add_14_36_groupi_n_2137), .y(csa_tree_add_14_36_groupi_n_1058));
xor2 csa_tree_add_14_36_groupi_g51974__1786 (.a(csa_tree_add_14_36_groupi_n_228), .b(csa_tree_add_14_36_groupi_n_2136), .y(csa_tree_add_14_36_groupi_n_1089));
xor2 csa_tree_add_14_36_groupi_g51975__5953 (.a(csa_tree_add_14_36_groupi_n_2143), .b(csa_tree_add_14_36_groupi_n_2149), .y(csa_tree_add_14_36_groupi_n_1057));
xor2 csa_tree_add_14_36_groupi_g51976__5703 (.a(csa_tree_add_14_36_groupi_n_2039), .b(csa_tree_add_14_36_groupi_n_2059), .y(csa_tree_add_14_36_groupi_n_1056));
xor2 csa_tree_add_14_36_groupi_g51977__7114 (.a(csa_tree_add_14_36_groupi_n_2078), .b(csa_tree_add_14_36_groupi_n_2103), .y(csa_tree_add_14_36_groupi_n_1055));
xor2 csa_tree_add_14_36_groupi_g51978__5266 (.a(csa_tree_add_14_36_groupi_n_2102), .b(csa_tree_add_14_36_groupi_n_2094), .y(csa_tree_add_14_36_groupi_n_1054));
xor2 csa_tree_add_14_36_groupi_g51979__2250 (.a(csa_tree_add_14_36_groupi_n_135), .b(csa_tree_add_14_36_groupi_n_2040), .y(csa_tree_add_14_36_groupi_n_2285));
xor2 csa_tree_add_14_36_groupi_g51980__6083 (.a(csa_tree_add_14_36_groupi_n_2069), .b(csa_tree_add_14_36_groupi_n_2063), .y(csa_tree_add_14_36_groupi_n_1053));
xor2 csa_tree_add_14_36_groupi_g51981__2703 (.a(csa_tree_add_14_36_groupi_n_897), .b(csa_tree_add_14_36_groupi_n_2062), .y(csa_tree_add_14_36_groupi_n_1088));
xor2 csa_tree_add_14_36_groupi_g51982__5795 (.a(csa_tree_add_14_36_groupi_n_2068), .b(csa_tree_add_14_36_groupi_n_2057), .y(csa_tree_add_14_36_groupi_n_1052));
xor2 csa_tree_add_14_36_groupi_g51983__7344 (.a(csa_tree_add_14_36_groupi_n_2076), .b(csa_tree_add_14_36_groupi_n_2134), .y(csa_tree_add_14_36_groupi_n_1051));
xor2 csa_tree_add_14_36_groupi_g51984__1840 (.a(csa_tree_add_14_36_groupi_n_2084), .b(csa_tree_add_14_36_groupi_n_2060), .y(csa_tree_add_14_36_groupi_n_1050));
xor2 csa_tree_add_14_36_groupi_g51985__5019 (.a(csa_tree_add_14_36_groupi_n_2116), .b(csa_tree_add_14_36_groupi_n_2054), .y(csa_tree_add_14_36_groupi_n_1049));
xor2 csa_tree_add_14_36_groupi_g51986__1857 (.a(csa_tree_add_14_36_groupi_n_2080), .b(csa_tree_add_14_36_groupi_n_2025), .y(csa_tree_add_14_36_groupi_n_1048));
xor2 csa_tree_add_14_36_groupi_g51987__9906 (.a(csa_tree_add_14_36_groupi_n_2082), .b(csa_tree_add_14_36_groupi_n_2024), .y(csa_tree_add_14_36_groupi_n_1047));
xor2 csa_tree_add_14_36_groupi_g51988__8780 (.a(csa_tree_add_14_36_groupi_n_2085), .b(csa_tree_add_14_36_groupi_n_2023), .y(csa_tree_add_14_36_groupi_n_1046));
xor2 csa_tree_add_14_36_groupi_g51989__4296 (.a(csa_tree_add_14_36_groupi_n_830), .b(csa_tree_add_14_36_groupi_n_900), .y(csa_tree_add_14_36_groupi_n_1087));
xor2 csa_tree_add_14_36_groupi_g51990__3772 (.a(csa_tree_add_14_36_groupi_n_137), .b(csa_tree_add_14_36_groupi_n_2075), .y(csa_tree_add_14_36_groupi_n_1086));
xor2 csa_tree_add_14_36_groupi_g51991__1474 (.a(csa_tree_add_14_36_groupi_n_504), .b(csa_tree_add_14_36_groupi_n_2032), .y(csa_tree_add_14_36_groupi_n_1085));
xor2 csa_tree_add_14_36_groupi_g51992__4547 (.a(csa_tree_add_14_36_groupi_n_507), .b(csa_tree_add_14_36_groupi_n_2071), .y(csa_tree_add_14_36_groupi_n_1084));
xor2 csa_tree_add_14_36_groupi_g51993__9682 (.a(csa_tree_add_14_36_groupi_n_502), .b(csa_tree_add_14_36_groupi_n_2074), .y(csa_tree_add_14_36_groupi_n_1083));
xor2 csa_tree_add_14_36_groupi_g51994__2683 (.a(csa_tree_add_14_36_groupi_n_818), .b(csa_tree_add_14_36_groupi_n_2049), .y(csa_tree_add_14_36_groupi_n_1082));
xor2 csa_tree_add_14_36_groupi_g51995__1309 (.a(csa_tree_add_14_36_groupi_n_41), .b(csa_tree_add_14_36_groupi_n_2081), .y(csa_tree_add_14_36_groupi_n_1081));
xor2 csa_tree_add_14_36_groupi_g51997__2900 (.a(csa_tree_add_14_36_groupi_n_227), .b(csa_tree_add_14_36_groupi_n_2043), .y(csa_tree_add_14_36_groupi_n_1080));
xor2 csa_tree_add_14_36_groupi_g51998__2391 (.a(csa_tree_add_14_36_groupi_n_817), .b(csa_tree_add_14_36_groupi_n_2055), .y(csa_tree_add_14_36_groupi_n_1079));
xor2 csa_tree_add_14_36_groupi_g51999__7675 (.a(csa_tree_add_14_36_groupi_n_506), .b(csa_tree_add_14_36_groupi_n_2041), .y(csa_tree_add_14_36_groupi_n_1078));
xor2 csa_tree_add_14_36_groupi_g52000__7118 (.a(csa_tree_add_14_36_groupi_n_505), .b(csa_tree_add_14_36_groupi_n_2087), .y(csa_tree_add_14_36_groupi_n_1077));
nand2 csa_tree_add_14_36_groupi_g52001__8757 (.a(csa_tree_add_14_36_groupi_n_935), .b(csa_tree_add_14_36_groupi_n_829), .y(csa_tree_add_14_36_groupi_n_1076));
xor2 csa_tree_add_14_36_groupi_g52002__1786 (.a(csa_tree_add_14_36_groupi_n_138), .b(csa_tree_add_14_36_groupi_n_2047), .y(csa_tree_add_14_36_groupi_n_1075));
inv csa_tree_add_14_36_groupi_g52003 (.a(csa_tree_add_14_36_groupi_n_1014), .y(csa_tree_add_14_36_groupi_n_1045));
inv csa_tree_add_14_36_groupi_g52004 (.a(csa_tree_add_14_36_groupi_n_1008), .y(csa_tree_add_14_36_groupi_n_1044));
inv csa_tree_add_14_36_groupi_g52005 (.a(csa_tree_add_14_36_groupi_n_1005), .y(csa_tree_add_14_36_groupi_n_1043));
inv csa_tree_add_14_36_groupi_g52006 (.a(csa_tree_add_14_36_groupi_n_1003), .y(csa_tree_add_14_36_groupi_n_1042));
inv csa_tree_add_14_36_groupi_g52007 (.a(csa_tree_add_14_36_groupi_n_1001), .y(csa_tree_add_14_36_groupi_n_1041));
inv csa_tree_add_14_36_groupi_g52008 (.a(csa_tree_add_14_36_groupi_n_1000), .y(csa_tree_add_14_36_groupi_n_1040));
inv csa_tree_add_14_36_groupi_g52009 (.a(csa_tree_add_14_36_groupi_n_996), .y(csa_tree_add_14_36_groupi_n_1039));
inv csa_tree_add_14_36_groupi_g52010 (.a(csa_tree_add_14_36_groupi_n_995), .y(csa_tree_add_14_36_groupi_n_1038));
inv csa_tree_add_14_36_groupi_g52011 (.a(csa_tree_add_14_36_groupi_n_989), .y(csa_tree_add_14_36_groupi_n_1037));
inv csa_tree_add_14_36_groupi_g52012 (.a(csa_tree_add_14_36_groupi_n_988), .y(csa_tree_add_14_36_groupi_n_1036));
inv csa_tree_add_14_36_groupi_g52014 (.a(csa_tree_add_14_36_groupi_n_985), .y(csa_tree_add_14_36_groupi_n_1034));
inv csa_tree_add_14_36_groupi_g52016 (.a(csa_tree_add_14_36_groupi_n_973), .y(csa_tree_add_14_36_groupi_n_1032));
inv csa_tree_add_14_36_groupi_g52017 (.a(csa_tree_add_14_36_groupi_n_1029), .y(csa_tree_add_14_36_groupi_n_1030));
inv csa_tree_add_14_36_groupi_g52018 (.a(csa_tree_add_14_36_groupi_n_1024), .y(csa_tree_add_14_36_groupi_n_1025));
inv csa_tree_add_14_36_groupi_g52019 (.a(csa_tree_add_14_36_groupi_n_1022), .y(csa_tree_add_14_36_groupi_n_1021));
nand2 csa_tree_add_14_36_groupi_g52020__5953 (.a(csa_tree_add_14_36_groupi_n_2068), .b(csa_tree_add_14_36_groupi_n_2057), .y(csa_tree_add_14_36_groupi_n_1020));
nand2 csa_tree_add_14_36_groupi_g52022__7114 (.a(csa_tree_add_14_36_groupi_n_2084), .b(csa_tree_add_14_36_groupi_n_2060), .y(csa_tree_add_14_36_groupi_n_1018));
nand2 csa_tree_add_14_36_groupi_g52023__5266 (.a(csa_tree_add_14_36_groupi_n_2035), .b(csa_tree_add_14_36_groupi_n_894), .y(csa_tree_add_14_36_groupi_n_1017));
nand2 csa_tree_add_14_36_groupi_g52024__2250 (.a(csa_tree_add_14_36_groupi_n_2072), .b(csa_tree_add_14_36_groupi_n_2050), .y(csa_tree_add_14_36_groupi_n_1016));
nand2 csa_tree_add_14_36_groupi_g52025__6083 (.a(csa_tree_add_14_36_groupi_n_2070), .b(csa_tree_add_14_36_groupi_n_2052), .y(csa_tree_add_14_36_groupi_n_1015));
nor2 csa_tree_add_14_36_groupi_g52026__2703 (.a(csa_tree_add_14_36_groupi_n_2083), .b(csa_tree_add_14_36_groupi_n_2137), .y(csa_tree_add_14_36_groupi_n_1014));
nand2 csa_tree_add_14_36_groupi_g52027__5795 (.a(csa_tree_add_14_36_groupi_n_2116), .b(csa_tree_add_14_36_groupi_n_2054), .y(csa_tree_add_14_36_groupi_n_1013));
nand2 csa_tree_add_14_36_groupi_g52028__7344 (.a(csa_tree_add_14_36_groupi_n_2078), .b(csa_tree_add_14_36_groupi_n_2103), .y(csa_tree_add_14_36_groupi_n_1012));
nor2 csa_tree_add_14_36_groupi_g52030__5019 (.a(csa_tree_add_14_36_groupi_n_261), .b(csa_tree_add_14_36_groupi_n_2032), .y(csa_tree_add_14_36_groupi_n_1010));
nand2 csa_tree_add_14_36_groupi_g52031__1857 (.a(csa_tree_add_14_36_groupi_n_2083), .b(csa_tree_add_14_36_groupi_n_2137), .y(csa_tree_add_14_36_groupi_n_1009));
nor2 csa_tree_add_14_36_groupi_g52032__9906 (.a(n_133), .b(csa_tree_add_14_36_groupi_n_2136), .y(csa_tree_add_14_36_groupi_n_1008));
nand2 csa_tree_add_14_36_groupi_g52033__8780 (.a(n_133), .b(csa_tree_add_14_36_groupi_n_2136), .y(csa_tree_add_14_36_groupi_n_1007));
nand2 csa_tree_add_14_36_groupi_g52034__4296 (.a(csa_tree_add_14_36_groupi_n_2038), .b(csa_tree_add_14_36_groupi_n_2045), .y(csa_tree_add_14_36_groupi_n_1006));
nor2 csa_tree_add_14_36_groupi_g52035__3772 (.a(csa_tree_add_14_36_groupi_n_2038), .b(csa_tree_add_14_36_groupi_n_2045), .y(csa_tree_add_14_36_groupi_n_1005));
nor2 csa_tree_add_14_36_groupi_g52037__4547 (.a(csa_tree_add_14_36_groupi_n_2072), .b(csa_tree_add_14_36_groupi_n_2050), .y(csa_tree_add_14_36_groupi_n_1003));
nand2 csa_tree_add_14_36_groupi_g52038__9682 (.a(csa_tree_add_14_36_groupi_n_2102), .b(csa_tree_add_14_36_groupi_n_2094), .y(csa_tree_add_14_36_groupi_n_1002));
nor2 csa_tree_add_14_36_groupi_g52039__2683 (.a(n_131), .b(csa_tree_add_14_36_groupi_n_2075), .y(csa_tree_add_14_36_groupi_n_1001));
nor2 csa_tree_add_14_36_groupi_g52040__1309 (.a(csa_tree_add_14_36_groupi_n_2085), .b(csa_tree_add_14_36_groupi_n_2023), .y(csa_tree_add_14_36_groupi_n_1000));
nor2 csa_tree_add_14_36_groupi_g52041__6877 (.a(csa_tree_add_14_36_groupi_n_2069), .b(csa_tree_add_14_36_groupi_n_2063), .y(csa_tree_add_14_36_groupi_n_999));
nand2 csa_tree_add_14_36_groupi_g52042__2900 (.a(csa_tree_add_14_36_groupi_n_2069), .b(csa_tree_add_14_36_groupi_n_2063), .y(csa_tree_add_14_36_groupi_n_998));
nand2 csa_tree_add_14_36_groupi_g52043__2391 (.a(n_129), .b(csa_tree_add_14_36_groupi_n_2047), .y(csa_tree_add_14_36_groupi_n_997));
nor2 csa_tree_add_14_36_groupi_g52044__7675 (.a(n_129), .b(csa_tree_add_14_36_groupi_n_2047), .y(csa_tree_add_14_36_groupi_n_996));
nor2 csa_tree_add_14_36_groupi_g52045__7118 (.a(csa_tree_add_14_36_groupi_n_2080), .b(csa_tree_add_14_36_groupi_n_2025), .y(csa_tree_add_14_36_groupi_n_995));
nand2 csa_tree_add_14_36_groupi_g52046__8757 (.a(csa_tree_add_14_36_groupi_n_2082), .b(csa_tree_add_14_36_groupi_n_2024), .y(csa_tree_add_14_36_groupi_n_994));
nor2 csa_tree_add_14_36_groupi_g52047__1786 (.a(csa_tree_add_14_36_groupi_n_2082), .b(csa_tree_add_14_36_groupi_n_2024), .y(csa_tree_add_14_36_groupi_n_993));
nor2 csa_tree_add_14_36_groupi_g52048__5953 (.a(csa_tree_add_14_36_groupi_n_2076), .b(csa_tree_add_14_36_groupi_n_2134), .y(csa_tree_add_14_36_groupi_n_992));
nand2 csa_tree_add_14_36_groupi_g52049__5703 (.a(csa_tree_add_14_36_groupi_n_2080), .b(csa_tree_add_14_36_groupi_n_2025), .y(csa_tree_add_14_36_groupi_n_991));
nand2 csa_tree_add_14_36_groupi_g52050__7114 (.a(csa_tree_add_14_36_groupi_n_2073), .b(csa_tree_add_14_36_groupi_n_2062), .y(csa_tree_add_14_36_groupi_n_990));
nor2 csa_tree_add_14_36_groupi_g52051__5266 (.a(csa_tree_add_14_36_groupi_n_2070), .b(csa_tree_add_14_36_groupi_n_2052), .y(csa_tree_add_14_36_groupi_n_989));
nor2 csa_tree_add_14_36_groupi_g52052__2250 (.a(csa_tree_add_14_36_groupi_n_2068), .b(csa_tree_add_14_36_groupi_n_2057), .y(csa_tree_add_14_36_groupi_n_988));
nand2 csa_tree_add_14_36_groupi_g52054__2703 (.a(csa_tree_add_14_36_groupi_n_2143), .b(csa_tree_add_14_36_groupi_n_2149), .y(csa_tree_add_14_36_groupi_n_986));
nor2 csa_tree_add_14_36_groupi_g52055__5795 (.a(csa_tree_add_14_36_groupi_n_2143), .b(csa_tree_add_14_36_groupi_n_2149), .y(csa_tree_add_14_36_groupi_n_985));
nor2 csa_tree_add_14_36_groupi_g52056__7344 (.a(csa_tree_add_14_36_groupi_n_2084), .b(csa_tree_add_14_36_groupi_n_2060), .y(csa_tree_add_14_36_groupi_n_984));
nor2 csa_tree_add_14_36_groupi_g52057__1840 (.a(csa_tree_add_14_36_groupi_n_2078), .b(csa_tree_add_14_36_groupi_n_2103), .y(csa_tree_add_14_36_groupi_n_983));
nand2 csa_tree_add_14_36_groupi_g52059__1857 (.a(csa_tree_add_14_36_groupi_n_2076), .b(csa_tree_add_14_36_groupi_n_2134), .y(csa_tree_add_14_36_groupi_n_981));
nand2 csa_tree_add_14_36_groupi_g52060__9906 (.a(csa_tree_add_14_36_groupi_n_2140), .b(csa_tree_add_14_36_groupi_n_2092), .y(csa_tree_add_14_36_groupi_n_980));
nand2 csa_tree_add_14_36_groupi_g52061__8780 (.a(csa_tree_add_14_36_groupi_n_2039), .b(csa_tree_add_14_36_groupi_n_2059), .y(csa_tree_add_14_36_groupi_n_979));
nand2 csa_tree_add_14_36_groupi_g52064__1474 (.a(n_131), .b(csa_tree_add_14_36_groupi_n_2075), .y(csa_tree_add_14_36_groupi_n_976));
nand2 csa_tree_add_14_36_groupi_g52065__4547 (.a(csa_tree_add_14_36_groupi_n_2085), .b(csa_tree_add_14_36_groupi_n_2023), .y(csa_tree_add_14_36_groupi_n_975));
nand2 csa_tree_add_14_36_groupi_g52066__9682 (.a(n_141), .b(csa_tree_add_14_36_groupi_n_2040), .y(csa_tree_add_14_36_groupi_n_974));
nor2 csa_tree_add_14_36_groupi_g52067__2683 (.a(n_141), .b(csa_tree_add_14_36_groupi_n_2040), .y(csa_tree_add_14_36_groupi_n_973));
nand2 csa_tree_add_14_36_groupi_g52068__1309 (.a(csa_tree_add_14_36_groupi_n_812), .b(csa_tree_add_14_36_groupi_n_2056), .y(csa_tree_add_14_36_groupi_n_972));
nor2 csa_tree_add_14_36_groupi_g52070__2900 (.a(csa_tree_add_14_36_groupi_n_262), .b(csa_tree_add_14_36_groupi_n_2041), .y(csa_tree_add_14_36_groupi_n_970));
nor2 csa_tree_add_14_36_groupi_g52071__2391 (.a(csa_tree_add_14_36_groupi_n_2034), .b(csa_tree_add_14_36_groupi_n_898), .y(csa_tree_add_14_36_groupi_n_969));
nand2 csa_tree_add_14_36_groupi_g52072__7675 (.a(csa_tree_add_14_36_groupi_n_413), .b(csa_tree_add_14_36_groupi_n_2071), .y(csa_tree_add_14_36_groupi_n_968));
nand2 csa_tree_add_14_36_groupi_g52073__7118 (.a(csa_tree_add_14_36_groupi_n_2033), .b(csa_tree_add_14_36_groupi_n_902), .y(csa_tree_add_14_36_groupi_n_1031));
nor2 csa_tree_add_14_36_groupi_g52074__8757 (.a(csa_tree_add_14_36_groupi_n_2029), .b(csa_tree_add_14_36_groupi_n_2053), .y(csa_tree_add_14_36_groupi_n_1029));
nand2 csa_tree_add_14_36_groupi_g52075__1786 (.a(csa_tree_add_14_36_groupi_n_803), .b(csa_tree_add_14_36_groupi_n_878), .y(csa_tree_add_14_36_groupi_n_1028));
nand2 csa_tree_add_14_36_groupi_g52076__5953 (.a(csa_tree_add_14_36_groupi_n_298), .b(csa_tree_add_14_36_groupi_n_2089), .y(csa_tree_add_14_36_groupi_n_1027));
nand2 csa_tree_add_14_36_groupi_g52077__5703 (.a(csa_tree_add_14_36_groupi_n_62), .b(csa_tree_add_14_36_groupi_n_2110), .y(csa_tree_add_14_36_groupi_n_1026));
nand2 csa_tree_add_14_36_groupi_g52078__7114 (.a(csa_tree_add_14_36_groupi_n_867), .b(csa_tree_add_14_36_groupi_n_748), .y(csa_tree_add_14_36_groupi_n_1024));
nand2 csa_tree_add_14_36_groupi_g52079__5266 (.a(csa_tree_add_14_36_groupi_n_866), .b(csa_tree_add_14_36_groupi_n_810), .y(csa_tree_add_14_36_groupi_n_1023));
nand2 csa_tree_add_14_36_groupi_g52080__2250 (.a(csa_tree_add_14_36_groupi_n_2029), .b(csa_tree_add_14_36_groupi_n_2053), .y(csa_tree_add_14_36_groupi_n_1022));
inv csa_tree_add_14_36_groupi_g52081 (.a(csa_tree_add_14_36_groupi_n_948), .y(csa_tree_add_14_36_groupi_n_967));
nand2 csa_tree_add_14_36_groupi_g52082__6083 (.a(csa_tree_add_14_36_groupi_n_749), .b(csa_tree_add_14_36_groupi_n_900), .y(csa_tree_add_14_36_groupi_n_962));
nand2 csa_tree_add_14_36_groupi_g52083__2703 (.a(csa_tree_add_14_36_groupi_n_799), .b(csa_tree_add_14_36_groupi_n_2055), .y(csa_tree_add_14_36_groupi_n_961));
nor2 csa_tree_add_14_36_groupi_g52084__5795 (.a(csa_tree_add_14_36_groupi_n_2155), .b(csa_tree_add_14_36_groupi_n_896), .y(csa_tree_add_14_36_groupi_n_960));
nand2 csa_tree_add_14_36_groupi_g52085__7344 (.a(csa_tree_add_14_36_groupi_n_750), .b(csa_tree_add_14_36_groupi_n_2049), .y(csa_tree_add_14_36_groupi_n_959));
nand2 csa_tree_add_14_36_groupi_g52086__1840 (.a(csa_tree_add_14_36_groupi_n_801), .b(csa_tree_add_14_36_groupi_n_889), .y(csa_tree_add_14_36_groupi_n_958));
nand2 csa_tree_add_14_36_groupi_g52087__5019 (.a(csa_tree_add_14_36_groupi_n_260), .b(csa_tree_add_14_36_groupi_n_2074), .y(csa_tree_add_14_36_groupi_n_957));
nor2 csa_tree_add_14_36_groupi_g52088__1857 (.a(csa_tree_add_14_36_groupi_n_2158), .b(csa_tree_add_14_36_groupi_n_895), .y(csa_tree_add_14_36_groupi_n_956));
nor2 csa_tree_add_14_36_groupi_g52089__9906 (.a(csa_tree_add_14_36_groupi_n_263), .b(csa_tree_add_14_36_groupi_n_2087), .y(csa_tree_add_14_36_groupi_n_955));
nand2 csa_tree_add_14_36_groupi_g52090__8780 (.a(csa_tree_add_14_36_groupi_n_868), .b(csa_tree_add_14_36_groupi_n_886), .y(csa_tree_add_14_36_groupi_n_954));
nand2 csa_tree_add_14_36_groupi_g52091__4296 (.a(csa_tree_add_14_36_groupi_n_726), .b(csa_tree_add_14_36_groupi_n_890), .y(csa_tree_add_14_36_groupi_n_953));
nor2 csa_tree_add_14_36_groupi_g52092__3772 (.a(csa_tree_add_14_36_groupi_n_863), .b(csa_tree_add_14_36_groupi_n_796), .y(csa_tree_add_14_36_groupi_n_952));
nand2 csa_tree_add_14_36_groupi_g52093__1474 (.a(csa_tree_add_14_36_groupi_n_860), .b(csa_tree_add_14_36_groupi_n_315), .y(csa_tree_add_14_36_groupi_n_951));
nand2 csa_tree_add_14_36_groupi_g52094__4547 (.a(csa_tree_add_14_36_groupi_n_888), .b(csa_tree_add_14_36_groupi_n_732), .y(csa_tree_add_14_36_groupi_n_950));
nand2 csa_tree_add_14_36_groupi_g52095__9682 (.a(csa_tree_add_14_36_groupi_n_730), .b(csa_tree_add_14_36_groupi_n_887), .y(csa_tree_add_14_36_groupi_n_949));
nor2 csa_tree_add_14_36_groupi_g52096__2683 (.a(csa_tree_add_14_36_groupi_n_727), .b(csa_tree_add_14_36_groupi_n_854), .y(csa_tree_add_14_36_groupi_n_948));
nand2 csa_tree_add_14_36_groupi_g52097__1309 (.a(csa_tree_add_14_36_groupi_n_723), .b(csa_tree_add_14_36_groupi_n_884), .y(csa_tree_add_14_36_groupi_n_947));
nand2 csa_tree_add_14_36_groupi_g52098__6877 (.a(csa_tree_add_14_36_groupi_n_725), .b(csa_tree_add_14_36_groupi_n_883), .y(csa_tree_add_14_36_groupi_n_946));
nand2 csa_tree_add_14_36_groupi_g52099__2900 (.a(csa_tree_add_14_36_groupi_n_722), .b(csa_tree_add_14_36_groupi_n_882), .y(csa_tree_add_14_36_groupi_n_945));
nand2 csa_tree_add_14_36_groupi_g52100__2391 (.a(csa_tree_add_14_36_groupi_n_885), .b(csa_tree_add_14_36_groupi_n_724), .y(csa_tree_add_14_36_groupi_n_944));
nand2 csa_tree_add_14_36_groupi_g52101__7675 (.a(csa_tree_add_14_36_groupi_n_731), .b(csa_tree_add_14_36_groupi_n_881), .y(csa_tree_add_14_36_groupi_n_943));
nand2 csa_tree_add_14_36_groupi_g52102__7118 (.a(csa_tree_add_14_36_groupi_n_721), .b(csa_tree_add_14_36_groupi_n_880), .y(csa_tree_add_14_36_groupi_n_942));
nand2 csa_tree_add_14_36_groupi_g52103__8757 (.a(n_2764), .b(csa_tree_add_14_36_groupi_n_879), .y(csa_tree_add_14_36_groupi_n_941));
nor2 csa_tree_add_14_36_groupi_g52104__1786 (.a(csa_tree_add_14_36_groupi_n_875), .b(csa_tree_add_14_36_groupi_n_709), .y(csa_tree_add_14_36_groupi_n_940));
nand2 csa_tree_add_14_36_groupi_g52105__5953 (.a(csa_tree_add_14_36_groupi_n_877), .b(csa_tree_add_14_36_groupi_n_798), .y(csa_tree_add_14_36_groupi_n_939));
nand2 csa_tree_add_14_36_groupi_g52106__5703 (.a(csa_tree_add_14_36_groupi_n_876), .b(csa_tree_add_14_36_groupi_n_794), .y(csa_tree_add_14_36_groupi_n_938));
nand2 csa_tree_add_14_36_groupi_g52107__7114 (.a(csa_tree_add_14_36_groupi_n_822), .b(n_2517), .y(csa_tree_add_14_36_groupi_n_937));
nand2 csa_tree_add_14_36_groupi_g52108__5266 (.a(csa_tree_add_14_36_groupi_n_823), .b(n_2522), .y(csa_tree_add_14_36_groupi_n_936));
nand2 csa_tree_add_14_36_groupi_g52109__2250 (.a(csa_tree_add_14_36_groupi_n_819), .b(csa_tree_add_14_36_groupi_n_729), .y(csa_tree_add_14_36_groupi_n_935));
nand2 csa_tree_add_14_36_groupi_g52110__6083 (.a(csa_tree_add_14_36_groupi_n_827), .b(n_2509), .y(csa_tree_add_14_36_groupi_n_934));
nand2 csa_tree_add_14_36_groupi_g52111__2703 (.a(csa_tree_add_14_36_groupi_n_826), .b(n_2620), .y(csa_tree_add_14_36_groupi_n_933));
xor2 csa_tree_add_14_36_groupi_g52112__5795 (.a(csa_tree_add_14_36_groupi_n_802), .b(csa_tree_add_14_36_groupi_n_316), .y(csa_tree_add_14_36_groupi_n_932));
nand2 csa_tree_add_14_36_groupi_g52113__7344 (.a(n_147), .b(csa_tree_add_14_36_groupi_n_904), .y(csa_tree_add_14_36_groupi_n_966));
xor2 csa_tree_add_14_36_groupi_g52114__1840 (.a(csa_tree_add_14_36_groupi_n_806), .b(csa_tree_add_14_36_groupi_n_103), .y(csa_tree_add_14_36_groupi_n_931));
nand2 csa_tree_add_14_36_groupi_g52115__5019 (.a(csa_tree_add_14_36_groupi_n_80), .b(csa_tree_add_14_36_groupi_n_2044), .y(csa_tree_add_14_36_groupi_n_930));
nand2 csa_tree_add_14_36_groupi_g52116__1857 (.a(csa_tree_add_14_36_groupi_n_892), .b(n_2698), .y(csa_tree_add_14_36_groupi_n_965));
nand2 csa_tree_add_14_36_groupi_g52122__4547 (.a(n_125), .b(csa_tree_add_14_36_groupi_n_901), .y(csa_tree_add_14_36_groupi_n_924));
xor2 csa_tree_add_14_36_groupi_g52123__9682 (.a(csa_tree_add_14_36_groupi_n_710), .b(csa_tree_add_14_36_groupi_n_777), .y(csa_tree_add_14_36_groupi_n_923));
xor2 csa_tree_add_14_36_groupi_g52124__2683 (.a(csa_tree_add_14_36_groupi_n_719), .b(csa_tree_add_14_36_groupi_n_794), .y(csa_tree_add_14_36_groupi_n_922));
xor2 csa_tree_add_14_36_groupi_g52125__1309 (.a(csa_tree_add_14_36_groupi_n_736), .b(csa_tree_add_14_36_groupi_n_709), .y(csa_tree_add_14_36_groupi_n_921));
xor2 csa_tree_add_14_36_groupi_g52126__6877 (.a(csa_tree_add_14_36_groupi_n_774), .b(csa_tree_add_14_36_groupi_n_775), .y(csa_tree_add_14_36_groupi_n_920));
xor2 csa_tree_add_14_36_groupi_g52127__2900 (.a(csa_tree_add_14_36_groupi_n_783), .b(csa_tree_add_14_36_groupi_n_702), .y(csa_tree_add_14_36_groupi_n_919));
xor2 csa_tree_add_14_36_groupi_g52128__2391 (.a(csa_tree_add_14_36_groupi_n_780), .b(csa_tree_add_14_36_groupi_n_705), .y(csa_tree_add_14_36_groupi_n_918));
xor2 csa_tree_add_14_36_groupi_g52129__7675 (.a(csa_tree_add_14_36_groupi_n_798), .b(csa_tree_add_14_36_groupi_n_703), .y(csa_tree_add_14_36_groupi_n_917));
xor2 csa_tree_add_14_36_groupi_g52130__7118 (.a(csa_tree_add_14_36_groupi_n_789), .b(csa_tree_add_14_36_groupi_n_712), .y(csa_tree_add_14_36_groupi_n_916));
xor2 csa_tree_add_14_36_groupi_g52131__8757 (.a(csa_tree_add_14_36_groupi_n_792), .b(csa_tree_add_14_36_groupi_n_704), .y(csa_tree_add_14_36_groupi_n_915));
xor2 csa_tree_add_14_36_groupi_g52133__5953 (.a(csa_tree_add_14_36_groupi_n_707), .b(csa_tree_add_14_36_groupi_n_706), .y(csa_tree_add_14_36_groupi_n_913));
xor2 csa_tree_add_14_36_groupi_g52134__5703 (.a(csa_tree_add_14_36_groupi_n_708), .b(csa_tree_add_14_36_groupi_n_650), .y(csa_tree_add_14_36_groupi_n_912));
xor2 csa_tree_add_14_36_groupi_g52135__7114 (.a(csa_tree_add_14_36_groupi_n_717), .b(csa_tree_add_14_36_groupi_n_720), .y(csa_tree_add_14_36_groupi_n_911));
xor2 csa_tree_add_14_36_groupi_g52136__5266 (.a(csa_tree_add_14_36_groupi_n_791), .b(csa_tree_add_14_36_groupi_n_732), .y(csa_tree_add_14_36_groupi_n_910));
xor2 csa_tree_add_14_36_groupi_g52137__2250 (.a(csa_tree_add_14_36_groupi_n_724), .b(csa_tree_add_14_36_groupi_n_715), .y(csa_tree_add_14_36_groupi_n_909));
xor2 csa_tree_add_14_36_groupi_g52138__6083 (.a(csa_tree_add_14_36_groupi_n_782), .b(csa_tree_add_14_36_groupi_n_716), .y(csa_tree_add_14_36_groupi_n_908));
xor2 csa_tree_add_14_36_groupi_g52139__2703 (.a(csa_tree_add_14_36_groupi_n_787), .b(csa_tree_add_14_36_groupi_n_651), .y(csa_tree_add_14_36_groupi_n_907));
xor2 csa_tree_add_14_36_groupi_g52140__5795 (.a(csa_tree_add_14_36_groupi_n_781), .b(csa_tree_add_14_36_groupi_n_786), .y(csa_tree_add_14_36_groupi_n_906));
xor2 csa_tree_add_14_36_groupi_g52141__7344 (.a(csa_tree_add_14_36_groupi_n_728), .b(csa_tree_add_14_36_groupi_n_2135), .y(csa_tree_add_14_36_groupi_n_905));
xor2 csa_tree_add_14_36_groupi_g52142__1840 (.a(n_79), .b(csa_tree_add_14_36_groupi_n_2106), .y(csa_tree_add_14_36_groupi_n_964));
xor2 csa_tree_add_14_36_groupi_g52143__5019 (.a(n_83), .b(csa_tree_add_14_36_groupi_n_2115), .y(csa_tree_add_14_36_groupi_n_963));
inv csa_tree_add_14_36_groupi_g52144 (.a(csa_tree_add_14_36_groupi_n_2110), .y(csa_tree_add_14_36_groupi_n_904));
inv csa_tree_add_14_36_groupi_g52145 (.a(csa_tree_add_14_36_groupi_n_2061), .y(csa_tree_add_14_36_groupi_n_903));
inv csa_tree_add_14_36_groupi_g52146 (.a(csa_tree_add_14_36_groupi_n_2089), .y(csa_tree_add_14_36_groupi_n_902));
inv csa_tree_add_14_36_groupi_g52147 (.a(csa_tree_add_14_36_groupi_n_2044), .y(csa_tree_add_14_36_groupi_n_901));
inv csa_tree_add_14_36_groupi_g52148 (.a(csa_tree_add_14_36_groupi_n_2032), .y(csa_tree_add_14_36_groupi_n_898));
inv csa_tree_add_14_36_groupi_g52149 (.a(csa_tree_add_14_36_groupi_n_2073), .y(csa_tree_add_14_36_groupi_n_897));
inv csa_tree_add_14_36_groupi_g52150 (.a(csa_tree_add_14_36_groupi_n_2041), .y(csa_tree_add_14_36_groupi_n_896));
inv csa_tree_add_14_36_groupi_g52151 (.a(csa_tree_add_14_36_groupi_n_2087), .y(csa_tree_add_14_36_groupi_n_895));
inv csa_tree_add_14_36_groupi_g52152 (.a(csa_tree_add_14_36_groupi_n_2074), .y(csa_tree_add_14_36_groupi_n_894));
nand2 csa_tree_add_14_36_groupi_g52154__9906 (.a(n_2696), .b(csa_tree_add_14_36_groupi_n_2086), .y(csa_tree_add_14_36_groupi_n_892));
nor2 csa_tree_add_14_36_groupi_g52155__8780 (.a(csa_tree_add_14_36_groupi_n_497), .b(csa_tree_add_14_36_groupi_n_784), .y(csa_tree_add_14_36_groupi_n_891));
nand2 csa_tree_add_14_36_groupi_g52164__4296 (.a(n_83), .b(csa_tree_add_14_36_groupi_n_2115), .y(csa_tree_add_14_36_groupi_n_900));
inv csa_tree_add_14_36_groupi_g52214 (.a(csa_tree_add_14_36_groupi_n_864), .y(csa_tree_add_14_36_groupi_n_890));
inv csa_tree_add_14_36_groupi_g52215 (.a(csa_tree_add_14_36_groupi_n_862), .y(csa_tree_add_14_36_groupi_n_889));
inv csa_tree_add_14_36_groupi_g52216 (.a(csa_tree_add_14_36_groupi_n_858), .y(csa_tree_add_14_36_groupi_n_888));
inv csa_tree_add_14_36_groupi_g52217 (.a(csa_tree_add_14_36_groupi_n_856), .y(csa_tree_add_14_36_groupi_n_887));
inv csa_tree_add_14_36_groupi_g52218 (.a(csa_tree_add_14_36_groupi_n_853), .y(csa_tree_add_14_36_groupi_n_886));
inv csa_tree_add_14_36_groupi_g52219 (.a(csa_tree_add_14_36_groupi_n_852), .y(csa_tree_add_14_36_groupi_n_885));
inv csa_tree_add_14_36_groupi_g52220 (.a(csa_tree_add_14_36_groupi_n_850), .y(csa_tree_add_14_36_groupi_n_884));
inv csa_tree_add_14_36_groupi_g52221 (.a(csa_tree_add_14_36_groupi_n_848), .y(csa_tree_add_14_36_groupi_n_883));
inv csa_tree_add_14_36_groupi_g52222 (.a(csa_tree_add_14_36_groupi_n_846), .y(csa_tree_add_14_36_groupi_n_882));
inv csa_tree_add_14_36_groupi_g52223 (.a(csa_tree_add_14_36_groupi_n_841), .y(csa_tree_add_14_36_groupi_n_881));
inv csa_tree_add_14_36_groupi_g52224 (.a(csa_tree_add_14_36_groupi_n_839), .y(csa_tree_add_14_36_groupi_n_880));
inv csa_tree_add_14_36_groupi_g52225 (.a(csa_tree_add_14_36_groupi_n_837), .y(csa_tree_add_14_36_groupi_n_879));
inv csa_tree_add_14_36_groupi_g52226 (.a(csa_tree_add_14_36_groupi_n_835), .y(csa_tree_add_14_36_groupi_n_878));
inv csa_tree_add_14_36_groupi_g52227 (.a(csa_tree_add_14_36_groupi_n_834), .y(csa_tree_add_14_36_groupi_n_877));
inv csa_tree_add_14_36_groupi_g52228 (.a(csa_tree_add_14_36_groupi_n_832), .y(csa_tree_add_14_36_groupi_n_876));
inv csa_tree_add_14_36_groupi_g52229 (.a(csa_tree_add_14_36_groupi_n_874), .y(csa_tree_add_14_36_groupi_n_875));
nand2 csa_tree_add_14_36_groupi_g52230__1474 (.a(csa_tree_add_14_36_groupi_n_753), .b(csa_tree_add_14_36_groupi_n_2079), .y(csa_tree_add_14_36_groupi_n_867));
nand2 csa_tree_add_14_36_groupi_g52231__4547 (.a(csa_tree_add_14_36_groupi_n_808), .b(csa_tree_add_14_36_groupi_n_2081), .y(csa_tree_add_14_36_groupi_n_866));
nand2 csa_tree_add_14_36_groupi_g52232__9682 (.a(csa_tree_add_14_36_groupi_n_708), .b(csa_tree_add_14_36_groupi_n_650), .y(csa_tree_add_14_36_groupi_n_865));
nor2 csa_tree_add_14_36_groupi_g52233__2683 (.a(csa_tree_add_14_36_groupi_n_708), .b(csa_tree_add_14_36_groupi_n_650), .y(csa_tree_add_14_36_groupi_n_864));
nor2 csa_tree_add_14_36_groupi_g52234__1309 (.a(n_2586), .b(csa_tree_add_14_36_groupi_n_618), .y(csa_tree_add_14_36_groupi_n_863));
nor2 csa_tree_add_14_36_groupi_g52235__6877 (.a(csa_tree_add_14_36_groupi_n_787), .b(csa_tree_add_14_36_groupi_n_651), .y(csa_tree_add_14_36_groupi_n_862));
nand2 csa_tree_add_14_36_groupi_g52236__2900 (.a(csa_tree_add_14_36_groupi_n_787), .b(csa_tree_add_14_36_groupi_n_651), .y(csa_tree_add_14_36_groupi_n_861));
nand2 csa_tree_add_14_36_groupi_g52237__2391 (.a(csa_tree_add_14_36_groupi_n_802), .b(csa_tree_add_14_36_groupi_n_239), .y(csa_tree_add_14_36_groupi_n_860));
nand2 csa_tree_add_14_36_groupi_g52238__7675 (.a(csa_tree_add_14_36_groupi_n_781), .b(csa_tree_add_14_36_groupi_n_786), .y(csa_tree_add_14_36_groupi_n_859));
nor2 csa_tree_add_14_36_groupi_g52239__7118 (.a(csa_tree_add_14_36_groupi_n_791), .b(csa_tree_add_14_36_groupi_n_785), .y(csa_tree_add_14_36_groupi_n_858));
nand2 csa_tree_add_14_36_groupi_g52240__8757 (.a(csa_tree_add_14_36_groupi_n_791), .b(csa_tree_add_14_36_groupi_n_785), .y(csa_tree_add_14_36_groupi_n_857));
nor2 csa_tree_add_14_36_groupi_g52241__1786 (.a(csa_tree_add_14_36_groupi_n_781), .b(csa_tree_add_14_36_groupi_n_786), .y(csa_tree_add_14_36_groupi_n_856));
nand2 csa_tree_add_14_36_groupi_g52242__5953 (.a(csa_tree_add_14_36_groupi_n_780), .b(csa_tree_add_14_36_groupi_n_705), .y(csa_tree_add_14_36_groupi_n_855));
nor2 csa_tree_add_14_36_groupi_g52243__5703 (.a(csa_tree_add_14_36_groupi_n_780), .b(csa_tree_add_14_36_groupi_n_705), .y(csa_tree_add_14_36_groupi_n_854));
nor2 csa_tree_add_14_36_groupi_g52244__7114 (.a(csa_tree_add_14_36_groupi_n_782), .b(csa_tree_add_14_36_groupi_n_716), .y(csa_tree_add_14_36_groupi_n_853));
nor2 csa_tree_add_14_36_groupi_g52245__5266 (.a(csa_tree_add_14_36_groupi_n_790), .b(csa_tree_add_14_36_groupi_n_715), .y(csa_tree_add_14_36_groupi_n_852));
nand2 csa_tree_add_14_36_groupi_g52246__2250 (.a(csa_tree_add_14_36_groupi_n_789), .b(csa_tree_add_14_36_groupi_n_712), .y(csa_tree_add_14_36_groupi_n_851));
nor2 csa_tree_add_14_36_groupi_g52247 (.a(csa_tree_add_14_36_groupi_n_789), .b(csa_tree_add_14_36_groupi_n_712), .y(csa_tree_add_14_36_groupi_n_850));
nand2 csa_tree_add_14_36_groupi_g52248 (.a(csa_tree_add_14_36_groupi_n_792), .b(csa_tree_add_14_36_groupi_n_704), .y(csa_tree_add_14_36_groupi_n_849));
nor2 csa_tree_add_14_36_groupi_g52249 (.a(csa_tree_add_14_36_groupi_n_792), .b(csa_tree_add_14_36_groupi_n_704), .y(csa_tree_add_14_36_groupi_n_848));
nand2 csa_tree_add_14_36_groupi_g52250 (.a(csa_tree_add_14_36_groupi_n_783), .b(csa_tree_add_14_36_groupi_n_702), .y(csa_tree_add_14_36_groupi_n_847));
nor2 csa_tree_add_14_36_groupi_g52251 (.a(csa_tree_add_14_36_groupi_n_783), .b(csa_tree_add_14_36_groupi_n_702), .y(csa_tree_add_14_36_groupi_n_846));
nand2 csa_tree_add_14_36_groupi_g52252 (.a(csa_tree_add_14_36_groupi_n_782), .b(csa_tree_add_14_36_groupi_n_716), .y(csa_tree_add_14_36_groupi_n_845));
nand2 csa_tree_add_14_36_groupi_g52253 (.a(csa_tree_add_14_36_groupi_n_790), .b(csa_tree_add_14_36_groupi_n_715), .y(csa_tree_add_14_36_groupi_n_844));
nand2 csa_tree_add_14_36_groupi_g52254 (.a(csa_tree_add_14_36_groupi_n_774), .b(csa_tree_add_14_36_groupi_n_775), .y(csa_tree_add_14_36_groupi_n_843));
nand2 csa_tree_add_14_36_groupi_g52255 (.a(csa_tree_add_14_36_groupi_n_707), .b(csa_tree_add_14_36_groupi_n_706), .y(csa_tree_add_14_36_groupi_n_842));
nor2 csa_tree_add_14_36_groupi_g52256 (.a(csa_tree_add_14_36_groupi_n_774), .b(csa_tree_add_14_36_groupi_n_775), .y(csa_tree_add_14_36_groupi_n_841));
nand2 csa_tree_add_14_36_groupi_g52257 (.a(csa_tree_add_14_36_groupi_n_703), .b(csa_tree_add_14_36_groupi_n_713), .y(csa_tree_add_14_36_groupi_n_840));
nor2 csa_tree_add_14_36_groupi_g52258 (.a(csa_tree_add_14_36_groupi_n_707), .b(csa_tree_add_14_36_groupi_n_706), .y(csa_tree_add_14_36_groupi_n_839));
nand2 csa_tree_add_14_36_groupi_g52259 (.a(csa_tree_add_14_36_groupi_n_714), .b(csa_tree_add_14_36_groupi_n_718), .y(csa_tree_add_14_36_groupi_n_838));
nor2 csa_tree_add_14_36_groupi_g52260 (.a(csa_tree_add_14_36_groupi_n_714), .b(csa_tree_add_14_36_groupi_n_718), .y(csa_tree_add_14_36_groupi_n_837));
nand2 csa_tree_add_14_36_groupi_g52261 (.a(csa_tree_add_14_36_groupi_n_711), .b(csa_tree_add_14_36_groupi_n_777), .y(csa_tree_add_14_36_groupi_n_836));
nor2 csa_tree_add_14_36_groupi_g52262 (.a(csa_tree_add_14_36_groupi_n_717), .b(csa_tree_add_14_36_groupi_n_720), .y(csa_tree_add_14_36_groupi_n_835));
nor2 csa_tree_add_14_36_groupi_g52263 (.a(csa_tree_add_14_36_groupi_n_703), .b(csa_tree_add_14_36_groupi_n_713), .y(csa_tree_add_14_36_groupi_n_834));
nor2 csa_tree_add_14_36_groupi_g52264 (.a(csa_tree_add_14_36_groupi_n_711), .b(csa_tree_add_14_36_groupi_n_777), .y(csa_tree_add_14_36_groupi_n_833));
nor2 csa_tree_add_14_36_groupi_g52265 (.a(csa_tree_add_14_36_groupi_n_719), .b(csa_tree_add_14_36_groupi_n_778), .y(csa_tree_add_14_36_groupi_n_832));
nand2 csa_tree_add_14_36_groupi_g52266 (.a(csa_tree_add_14_36_groupi_n_719), .b(csa_tree_add_14_36_groupi_n_778), .y(csa_tree_add_14_36_groupi_n_831));
xor2 csa_tree_add_14_36_groupi_g52267 (.a(n_82), .b(csa_tree_add_14_36_groupi_n_2157), .y(csa_tree_add_14_36_groupi_n_830));
nand2 csa_tree_add_14_36_groupi_g52268 (.a(csa_tree_add_14_36_groupi_n_806), .b(csa_tree_add_14_36_groupi_n_104), .y(csa_tree_add_14_36_groupi_n_829));
nand2 csa_tree_add_14_36_groupi_g52269 (.a(n_2507), .b(csa_tree_add_14_36_groupi_n_112), .y(csa_tree_add_14_36_groupi_n_828));
nand2 csa_tree_add_14_36_groupi_g52270 (.a(csa_tree_add_14_36_groupi_n_738), .b(n_2508), .y(csa_tree_add_14_36_groupi_n_827));
nand2 csa_tree_add_14_36_groupi_g52271 (.a(csa_tree_add_14_36_groupi_n_740), .b(csa_tree_add_14_36_groupi_n_101), .y(csa_tree_add_14_36_groupi_n_826));
nor2 csa_tree_add_14_36_groupi_g52272 (.a(csa_tree_add_14_36_groupi_n_743), .b(n_2526), .y(csa_tree_add_14_36_groupi_n_825));
nand2 csa_tree_add_14_36_groupi_g52273 (.a(n_2520), .b(csa_tree_add_14_36_groupi_n_107), .y(csa_tree_add_14_36_groupi_n_824));
nand2 csa_tree_add_14_36_groupi_g52274 (.a(csa_tree_add_14_36_groupi_n_744), .b(n_2521), .y(csa_tree_add_14_36_groupi_n_823));
nand2 csa_tree_add_14_36_groupi_g52275 (.a(csa_tree_add_14_36_groupi_n_746), .b(n_2516), .y(csa_tree_add_14_36_groupi_n_822));
nand2 csa_tree_add_14_36_groupi_g52276 (.a(csa_tree_add_14_36_groupi_n_741), .b(csa_tree_add_14_36_groupi_n_102), .y(csa_tree_add_14_36_groupi_n_821));
nand2 csa_tree_add_14_36_groupi_g52277 (.a(n_2515), .b(csa_tree_add_14_36_groupi_n_109), .y(csa_tree_add_14_36_groupi_n_820));
nand2 csa_tree_add_14_36_groupi_g52278 (.a(csa_tree_add_14_36_groupi_n_717), .b(csa_tree_add_14_36_groupi_n_720), .y(csa_tree_add_14_36_groupi_n_874));
nand2 csa_tree_add_14_36_groupi_g52279 (.a(csa_tree_add_14_36_groupi_n_805), .b(csa_tree_add_14_36_groupi_n_103), .y(csa_tree_add_14_36_groupi_n_819));
xor2 csa_tree_add_14_36_groupi_g52280 (.a(n_76), .b(csa_tree_add_14_36_groupi_n_2156), .y(csa_tree_add_14_36_groupi_n_818));
xor2 csa_tree_add_14_36_groupi_g52281 (.a(n_80), .b(csa_tree_add_14_36_groupi_n_2154), .y(csa_tree_add_14_36_groupi_n_817));
nand2 csa_tree_add_14_36_groupi_g52282 (.a(csa_tree_add_14_36_groupi_n_812), .b(csa_tree_add_14_36_groupi_n_813), .y(csa_tree_add_14_36_groupi_n_816));
xor2 csa_tree_add_14_36_groupi_g52284 (.a(csa_tree_add_14_36_groupi_n_83), .b(csa_tree_add_14_36_groupi_n_2026), .y(csa_tree_add_14_36_groupi_n_814));
xor2 csa_tree_add_14_36_groupi_g52286 (.a(n_159), .b(csa_tree_add_14_36_groupi_n_2065), .y(csa_tree_add_14_36_groupi_n_873));
xor2 csa_tree_add_14_36_groupi_g52287 (.a(n_81), .b(csa_tree_add_14_36_groupi_n_2051), .y(csa_tree_add_14_36_groupi_n_872));
xor2 csa_tree_add_14_36_groupi_g52288 (.a(n_157), .b(csa_tree_add_14_36_groupi_n_2124), .y(csa_tree_add_14_36_groupi_n_871));
xor2 csa_tree_add_14_36_groupi_g52289 (.a(n_77), .b(csa_tree_add_14_36_groupi_n_2123), .y(csa_tree_add_14_36_groupi_n_870));
xor2 csa_tree_add_14_36_groupi_g52290 (.a(n_155), .b(csa_tree_add_14_36_groupi_n_2030), .y(csa_tree_add_14_36_groupi_n_869));
nand2 csa_tree_add_14_36_groupi_g52291 (.a(csa_tree_add_14_36_groupi_n_693), .b(csa_tree_add_14_36_groupi_n_662), .y(csa_tree_add_14_36_groupi_n_868));
inv csa_tree_add_14_36_groupi_g52294 (.a(csa_tree_add_14_36_groupi_n_2077), .y(csa_tree_add_14_36_groupi_n_807));
inv csa_tree_add_14_36_groupi_g52295 (.a(csa_tree_add_14_36_groupi_n_806), .y(csa_tree_add_14_36_groupi_n_805));
inv csa_tree_add_14_36_groupi_g52296 (.a(csa_tree_add_14_36_groupi_n_799), .y(csa_tree_add_14_36_groupi_n_800));
inv csa_tree_add_14_36_groupi_g52297 (.a(n_2527), .y(csa_tree_add_14_36_groupi_n_796));
inv csa_tree_add_14_36_groupi_g52298 (.a(csa_tree_add_14_36_groupi_n_2135), .y(csa_tree_add_14_36_groupi_n_784));
nand2 csa_tree_add_14_36_groupi_g52300 (.a(csa_tree_add_14_36_groupi_n_577), .b(csa_tree_add_14_36_groupi_n_430), .y(csa_tree_add_14_36_groupi_n_771));
nand2 csa_tree_add_14_36_groupi_g52301 (.a(csa_tree_add_14_36_groupi_n_648), .b(csa_tree_add_14_36_groupi_n_385), .y(csa_tree_add_14_36_groupi_n_770));
nand2 csa_tree_add_14_36_groupi_g52302 (.a(csa_tree_add_14_36_groupi_n_560), .b(csa_tree_add_14_36_groupi_n_488), .y(csa_tree_add_14_36_groupi_n_769));
nand2 csa_tree_add_14_36_groupi_g52303 (.a(csa_tree_add_14_36_groupi_n_640), .b(csa_tree_add_14_36_groupi_n_431), .y(csa_tree_add_14_36_groupi_n_768));
nand2 csa_tree_add_14_36_groupi_g52304 (.a(csa_tree_add_14_36_groupi_n_639), .b(csa_tree_add_14_36_groupi_n_384), .y(csa_tree_add_14_36_groupi_n_767));
nand2 csa_tree_add_14_36_groupi_g52305 (.a(csa_tree_add_14_36_groupi_n_584), .b(csa_tree_add_14_36_groupi_n_451), .y(csa_tree_add_14_36_groupi_n_766));
nand2 csa_tree_add_14_36_groupi_g52306 (.a(csa_tree_add_14_36_groupi_n_585), .b(csa_tree_add_14_36_groupi_n_437), .y(csa_tree_add_14_36_groupi_n_765));
nand2 csa_tree_add_14_36_groupi_g52307 (.a(csa_tree_add_14_36_groupi_n_586), .b(csa_tree_add_14_36_groupi_n_461), .y(csa_tree_add_14_36_groupi_n_764));
nand2 csa_tree_add_14_36_groupi_g52308 (.a(csa_tree_add_14_36_groupi_n_587), .b(csa_tree_add_14_36_groupi_n_462), .y(csa_tree_add_14_36_groupi_n_763));
nand2 csa_tree_add_14_36_groupi_g52309 (.a(csa_tree_add_14_36_groupi_n_619), .b(csa_tree_add_14_36_groupi_n_442), .y(csa_tree_add_14_36_groupi_n_762));
nand2 csa_tree_add_14_36_groupi_g52310 (.a(csa_tree_add_14_36_groupi_n_594), .b(csa_tree_add_14_36_groupi_n_460), .y(csa_tree_add_14_36_groupi_n_761));
nand2 csa_tree_add_14_36_groupi_g52311 (.a(csa_tree_add_14_36_groupi_n_608), .b(csa_tree_add_14_36_groupi_n_443), .y(csa_tree_add_14_36_groupi_n_760));
nand2 csa_tree_add_14_36_groupi_g52312 (.a(csa_tree_add_14_36_groupi_n_610), .b(csa_tree_add_14_36_groupi_n_496), .y(csa_tree_add_14_36_groupi_n_759));
nand2 csa_tree_add_14_36_groupi_g52313 (.a(csa_tree_add_14_36_groupi_n_597), .b(csa_tree_add_14_36_groupi_n_440), .y(csa_tree_add_14_36_groupi_n_758));
nand2 csa_tree_add_14_36_groupi_g52314 (.a(csa_tree_add_14_36_groupi_n_649), .b(csa_tree_add_14_36_groupi_n_458), .y(csa_tree_add_14_36_groupi_n_757));
nand2 csa_tree_add_14_36_groupi_g52315 (.a(csa_tree_add_14_36_groupi_n_611), .b(csa_tree_add_14_36_groupi_n_455), .y(csa_tree_add_14_36_groupi_n_756));
nand2 csa_tree_add_14_36_groupi_g52316 (.a(csa_tree_add_14_36_groupi_n_609), .b(csa_tree_add_14_36_groupi_n_435), .y(csa_tree_add_14_36_groupi_n_755));
nand2 csa_tree_add_14_36_groupi_g52317 (.a(csa_tree_add_14_36_groupi_n_612), .b(csa_tree_add_14_36_groupi_n_463), .y(csa_tree_add_14_36_groupi_n_754));
nand2 csa_tree_add_14_36_groupi_g52318 (.a(n_78), .b(csa_tree_add_14_36_groupi_n_655), .y(csa_tree_add_14_36_groupi_n_813));
nand2 csa_tree_add_14_36_groupi_g52319 (.a(csa_tree_add_14_36_groupi_n_83), .b(csa_tree_add_14_36_groupi_n_2026), .y(csa_tree_add_14_36_groupi_n_753));
nand2 csa_tree_add_14_36_groupi_g52320 (.a(csa_tree_add_14_36_groupi_n_73), .b(csa_tree_add_14_36_groupi_n_2260), .y(csa_tree_add_14_36_groupi_n_812));
nand2 csa_tree_add_14_36_groupi_g52321 (.a(n_76), .b(csa_tree_add_14_36_groupi_n_657), .y(csa_tree_add_14_36_groupi_n_752));
nand2 csa_tree_add_14_36_groupi_g52323 (.a(n_121), .b(csa_tree_add_14_36_groupi_n_658), .y(csa_tree_add_14_36_groupi_n_810));
nand2 csa_tree_add_14_36_groupi_g52325 (.a(csa_tree_add_14_36_groupi_n_86), .b(csa_tree_add_14_36_groupi_n_2153), .y(csa_tree_add_14_36_groupi_n_808));
nand2 csa_tree_add_14_36_groupi_g52327 (.a(csa_tree_add_14_36_groupi_n_82), .b(csa_tree_add_14_36_groupi_n_2157), .y(csa_tree_add_14_36_groupi_n_751));
nand2 csa_tree_add_14_36_groupi_g52328 (.a(csa_tree_add_14_36_groupi_n_67), .b(csa_tree_add_14_36_groupi_n_2156), .y(csa_tree_add_14_36_groupi_n_750));
nand2 csa_tree_add_14_36_groupi_g52329 (.a(csa_tree_add_14_36_groupi_n_636), .b(csa_tree_add_14_36_groupi_n_614), .y(csa_tree_add_14_36_groupi_n_806));
nand2 csa_tree_add_14_36_groupi_g52330 (.a(n_82), .b(csa_tree_add_14_36_groupi_n_654), .y(csa_tree_add_14_36_groupi_n_749));
nand2 csa_tree_add_14_36_groupi_g52331 (.a(n_75), .b(csa_tree_add_14_36_groupi_n_661), .y(csa_tree_add_14_36_groupi_n_748));
nand2 csa_tree_add_14_36_groupi_g52333 (.a(csa_tree_add_14_36_groupi_n_617), .b(csa_tree_add_14_36_groupi_n_485), .y(csa_tree_add_14_36_groupi_n_2272));
nand2 csa_tree_add_14_36_groupi_g52336 (.a(csa_tree_add_14_36_groupi_n_635), .b(csa_tree_add_14_36_groupi_n_345), .y(csa_tree_add_14_36_groupi_n_803));
nand2 csa_tree_add_14_36_groupi_g52337 (.a(csa_tree_add_14_36_groupi_n_600), .b(csa_tree_add_14_36_groupi_n_459), .y(csa_tree_add_14_36_groupi_n_802));
nand2 csa_tree_add_14_36_groupi_g52338 (.a(csa_tree_add_14_36_groupi_n_637), .b(csa_tree_add_14_36_groupi_n_356), .y(csa_tree_add_14_36_groupi_n_801));
nand2 csa_tree_add_14_36_groupi_g52339 (.a(csa_tree_add_14_36_groupi_n_69), .b(csa_tree_add_14_36_groupi_n_2154), .y(csa_tree_add_14_36_groupi_n_799));
nand2 csa_tree_add_14_36_groupi_g52341 (.a(csa_tree_add_14_36_groupi_n_595), .b(csa_tree_add_14_36_groupi_n_456), .y(csa_tree_add_14_36_groupi_n_798));
nand2 csa_tree_add_14_36_groupi_g52346 (.a(csa_tree_add_14_36_groupi_n_541), .b(csa_tree_add_14_36_groupi_n_432), .y(csa_tree_add_14_36_groupi_n_794));
nand2 csa_tree_add_14_36_groupi_g52347 (.a(n_80), .b(csa_tree_add_14_36_groupi_n_653), .y(csa_tree_add_14_36_groupi_n_793));
nand2 csa_tree_add_14_36_groupi_g52348 (.a(csa_tree_add_14_36_groupi_n_591), .b(csa_tree_add_14_36_groupi_n_452), .y(csa_tree_add_14_36_groupi_n_792));
nand2 csa_tree_add_14_36_groupi_g52349 (.a(csa_tree_add_14_36_groupi_n_603), .b(csa_tree_add_14_36_groupi_n_444), .y(csa_tree_add_14_36_groupi_n_791));
nand2 csa_tree_add_14_36_groupi_g52350 (.a(csa_tree_add_14_36_groupi_n_606), .b(csa_tree_add_14_36_groupi_n_436), .y(csa_tree_add_14_36_groupi_n_790));
nand2 csa_tree_add_14_36_groupi_g52351 (.a(csa_tree_add_14_36_groupi_n_598), .b(csa_tree_add_14_36_groupi_n_447), .y(csa_tree_add_14_36_groupi_n_789));
nand2 csa_tree_add_14_36_groupi_g52352 (.a(n_155), .b(csa_tree_add_14_36_groupi_n_2030), .y(csa_tree_add_14_36_groupi_n_788));
nand2 csa_tree_add_14_36_groupi_g52353 (.a(csa_tree_add_14_36_groupi_n_604), .b(csa_tree_add_14_36_groupi_n_464), .y(csa_tree_add_14_36_groupi_n_787));
nand2 csa_tree_add_14_36_groupi_g52354 (.a(csa_tree_add_14_36_groupi_n_592), .b(csa_tree_add_14_36_groupi_n_439), .y(csa_tree_add_14_36_groupi_n_786));
nand2 csa_tree_add_14_36_groupi_g52355 (.a(csa_tree_add_14_36_groupi_n_602), .b(csa_tree_add_14_36_groupi_n_445), .y(csa_tree_add_14_36_groupi_n_785));
nand2 csa_tree_add_14_36_groupi_g52359 (.a(csa_tree_add_14_36_groupi_n_593), .b(csa_tree_add_14_36_groupi_n_441), .y(csa_tree_add_14_36_groupi_n_783));
nand2 csa_tree_add_14_36_groupi_g52360 (.a(csa_tree_add_14_36_groupi_n_599), .b(csa_tree_add_14_36_groupi_n_446), .y(csa_tree_add_14_36_groupi_n_782));
nand2 csa_tree_add_14_36_groupi_g52361 (.a(csa_tree_add_14_36_groupi_n_601), .b(csa_tree_add_14_36_groupi_n_438), .y(csa_tree_add_14_36_groupi_n_781));
nand2 csa_tree_add_14_36_groupi_g52366 (.a(csa_tree_add_14_36_groupi_n_590), .b(csa_tree_add_14_36_groupi_n_448), .y(csa_tree_add_14_36_groupi_n_780));
nand2 csa_tree_add_14_36_groupi_g52367 (.a(n_81), .b(csa_tree_add_14_36_groupi_n_660), .y(csa_tree_add_14_36_groupi_n_779));
nand2 csa_tree_add_14_36_groupi_g52368 (.a(csa_tree_add_14_36_groupi_n_605), .b(csa_tree_add_14_36_groupi_n_457), .y(csa_tree_add_14_36_groupi_n_778));
nand2 csa_tree_add_14_36_groupi_g52369 (.a(csa_tree_add_14_36_groupi_n_607), .b(csa_tree_add_14_36_groupi_n_453), .y(csa_tree_add_14_36_groupi_n_777));
nor2 csa_tree_add_14_36_groupi_g52370 (.a(csa_tree_add_14_36_groupi_n_70), .b(csa_tree_add_14_36_groupi_n_2065), .y(csa_tree_add_14_36_groupi_n_776));
nand2 csa_tree_add_14_36_groupi_g52371 (.a(csa_tree_add_14_36_groupi_n_644), .b(csa_tree_add_14_36_groupi_n_426), .y(csa_tree_add_14_36_groupi_n_775));
nand2 csa_tree_add_14_36_groupi_g52372 (.a(csa_tree_add_14_36_groupi_n_647), .b(csa_tree_add_14_36_groupi_n_429), .y(csa_tree_add_14_36_groupi_n_774));
inv csa_tree_add_14_36_groupi_g52377 (.a(n_2515), .y(csa_tree_add_14_36_groupi_n_746));
inv csa_tree_add_14_36_groupi_g52378 (.a(n_2520), .y(csa_tree_add_14_36_groupi_n_744));
inv csa_tree_add_14_36_groupi_g52379 (.a(n_2525), .y(csa_tree_add_14_36_groupi_n_743));
inv csa_tree_add_14_36_groupi_g52380 (.a(csa_tree_add_14_36_groupi_n_741), .y(csa_tree_add_14_36_groupi_n_740));
inv csa_tree_add_14_36_groupi_g52381 (.a(n_2507), .y(csa_tree_add_14_36_groupi_n_738));
inv csa_tree_add_14_36_groupi_g52382 (.a(csa_tree_add_14_36_groupi_n_711), .y(csa_tree_add_14_36_groupi_n_710));
nand2 csa_tree_add_14_36_groupi_g52383 (.a(csa_tree_add_14_36_groupi_n_538), .b(csa_tree_add_14_36_groupi_n_493), .y(csa_tree_add_14_36_groupi_n_701));
nand2 csa_tree_add_14_36_groupi_g52385 (.a(n_2461), .b(b_5), .y(csa_tree_add_14_36_groupi_n_699));
nand2 csa_tree_add_14_36_groupi_g52386 (.a(csa_tree_add_14_36_groupi_n_579), .b(csa_tree_add_14_36_groupi_n_393), .y(csa_tree_add_14_36_groupi_n_698));
nand2 csa_tree_add_14_36_groupi_g52387 (.a(csa_tree_add_14_36_groupi_n_537), .b(csa_tree_add_14_36_groupi_n_414), .y(csa_tree_add_14_36_groupi_n_697));
nand2 csa_tree_add_14_36_groupi_g52389 (.a(n_2675), .b(b_13), .y(csa_tree_add_14_36_groupi_n_695));
nand2 csa_tree_add_14_36_groupi_g52390 (.a(csa_tree_add_14_36_groupi_n_559), .b(csa_tree_add_14_36_groupi_n_392), .y(csa_tree_add_14_36_groupi_n_694));
nor2 csa_tree_add_14_36_groupi_g52391 (.a(csa_tree_add_14_36_groupi_n_518), .b(csa_tree_add_14_36_groupi_n_321), .y(csa_tree_add_14_36_groupi_n_693));
nand2 csa_tree_add_14_36_groupi_g52392 (.a(csa_tree_add_14_36_groupi_n_531), .b(csa_tree_add_14_36_groupi_n_357), .y(csa_tree_add_14_36_groupi_n_692));
nand2 csa_tree_add_14_36_groupi_g52394 (.a(csa_tree_add_14_36_groupi_n_516), .b(csa_tree_add_14_36_groupi_n_318), .y(csa_tree_add_14_36_groupi_n_690));
nand2 csa_tree_add_14_36_groupi_g52395 (.a(csa_tree_add_14_36_groupi_n_522), .b(csa_tree_add_14_36_groupi_n_337), .y(csa_tree_add_14_36_groupi_n_689));
nand2 csa_tree_add_14_36_groupi_g52396 (.a(csa_tree_add_14_36_groupi_n_638), .b(csa_tree_add_14_36_groupi_n_434), .y(csa_tree_add_14_36_groupi_n_688));
nand2 csa_tree_add_14_36_groupi_g52397 (.a(csa_tree_add_14_36_groupi_n_524), .b(csa_tree_add_14_36_groupi_n_408), .y(csa_tree_add_14_36_groupi_n_687));
nand2 csa_tree_add_14_36_groupi_g52398 (.a(csa_tree_add_14_36_groupi_n_525), .b(csa_tree_add_14_36_groupi_n_408), .y(csa_tree_add_14_36_groupi_n_686));
nand2 csa_tree_add_14_36_groupi_g52399 (.a(csa_tree_add_14_36_groupi_n_581), .b(csa_tree_add_14_36_groupi_n_425), .y(csa_tree_add_14_36_groupi_n_685));
nand2 csa_tree_add_14_36_groupi_g52400 (.a(csa_tree_add_14_36_groupi_n_544), .b(csa_tree_add_14_36_groupi_n_376), .y(csa_tree_add_14_36_groupi_n_684));
nand2 csa_tree_add_14_36_groupi_g52401 (.a(csa_tree_add_14_36_groupi_n_539), .b(csa_tree_add_14_36_groupi_n_380), .y(csa_tree_add_14_36_groupi_n_683));
nand2 csa_tree_add_14_36_groupi_g52402 (.a(csa_tree_add_14_36_groupi_n_570), .b(csa_tree_add_14_36_groupi_n_424), .y(csa_tree_add_14_36_groupi_n_682));
nand2 csa_tree_add_14_36_groupi_g52403 (.a(csa_tree_add_14_36_groupi_n_569), .b(csa_tree_add_14_36_groupi_n_375), .y(csa_tree_add_14_36_groupi_n_681));
nand2 csa_tree_add_14_36_groupi_g52404 (.a(csa_tree_add_14_36_groupi_n_536), .b(csa_tree_add_14_36_groupi_n_423), .y(csa_tree_add_14_36_groupi_n_680));
nand2 csa_tree_add_14_36_groupi_g52405 (.a(csa_tree_add_14_36_groupi_n_572), .b(csa_tree_add_14_36_groupi_n_374), .y(csa_tree_add_14_36_groupi_n_679));
nand2 csa_tree_add_14_36_groupi_g52406 (.a(csa_tree_add_14_36_groupi_n_534), .b(csa_tree_add_14_36_groupi_n_433), .y(csa_tree_add_14_36_groupi_n_678));
nand2 csa_tree_add_14_36_groupi_g52407 (.a(csa_tree_add_14_36_groupi_n_533), .b(csa_tree_add_14_36_groupi_n_389), .y(csa_tree_add_14_36_groupi_n_677));
nand2 csa_tree_add_14_36_groupi_g52408 (.a(csa_tree_add_14_36_groupi_n_540), .b(csa_tree_add_14_36_groupi_n_421), .y(csa_tree_add_14_36_groupi_n_676));
nand2 csa_tree_add_14_36_groupi_g52409 (.a(csa_tree_add_14_36_groupi_n_543), .b(csa_tree_add_14_36_groupi_n_379), .y(csa_tree_add_14_36_groupi_n_675));
nand2 csa_tree_add_14_36_groupi_g52410 (.a(csa_tree_add_14_36_groupi_n_645), .b(csa_tree_add_14_36_groupi_n_355), .y(csa_tree_add_14_36_groupi_n_674));
nand2 csa_tree_add_14_36_groupi_g52411 (.a(csa_tree_add_14_36_groupi_n_646), .b(csa_tree_add_14_36_groupi_n_340), .y(csa_tree_add_14_36_groupi_n_673));
nand2 csa_tree_add_14_36_groupi_g52412 (.a(csa_tree_add_14_36_groupi_n_558), .b(csa_tree_add_14_36_groupi_n_411), .y(csa_tree_add_14_36_groupi_n_672));
nand2 csa_tree_add_14_36_groupi_g52413 (.a(csa_tree_add_14_36_groupi_n_551), .b(csa_tree_add_14_36_groupi_n_343), .y(csa_tree_add_14_36_groupi_n_671));
nand2 csa_tree_add_14_36_groupi_g52414 (.a(csa_tree_add_14_36_groupi_n_550), .b(csa_tree_add_14_36_groupi_n_342), .y(csa_tree_add_14_36_groupi_n_670));
nand2 csa_tree_add_14_36_groupi_g52415 (.a(csa_tree_add_14_36_groupi_n_529), .b(csa_tree_add_14_36_groupi_n_338), .y(csa_tree_add_14_36_groupi_n_669));
nand2 csa_tree_add_14_36_groupi_g52416 (.a(csa_tree_add_14_36_groupi_n_589), .b(csa_tree_add_14_36_groupi_n_327), .y(csa_tree_add_14_36_groupi_n_668));
nand2 csa_tree_add_14_36_groupi_g52417 (.a(csa_tree_add_14_36_groupi_n_588), .b(csa_tree_add_14_36_groupi_n_328), .y(csa_tree_add_14_36_groupi_n_667));
nand2 csa_tree_add_14_36_groupi_g52418 (.a(csa_tree_add_14_36_groupi_n_643), .b(csa_tree_add_14_36_groupi_n_326), .y(csa_tree_add_14_36_groupi_n_666));
nand2 csa_tree_add_14_36_groupi_g52419 (.a(csa_tree_add_14_36_groupi_n_520), .b(csa_tree_add_14_36_groupi_n_335), .y(csa_tree_add_14_36_groupi_n_665));
nand2 csa_tree_add_14_36_groupi_g52420 (.a(csa_tree_add_14_36_groupi_n_532), .b(csa_tree_add_14_36_groupi_n_352), .y(csa_tree_add_14_36_groupi_n_664));
nand2 csa_tree_add_14_36_groupi_g52421 (.a(csa_tree_add_14_36_groupi_n_580), .b(csa_tree_add_14_36_groupi_n_418), .y(csa_tree_add_14_36_groupi_n_663));
nand2 csa_tree_add_14_36_groupi_g52425 (.a(csa_tree_add_14_36_groupi_n_517), .b(csa_tree_add_14_36_groupi_n_336), .y(csa_tree_add_14_36_groupi_n_741));
nand2 csa_tree_add_14_36_groupi_g52428 (.a(csa_tree_add_14_36_groupi_n_554), .b(csa_tree_add_14_36_groupi_n_353), .y(csa_tree_add_14_36_groupi_n_736));
nand2 csa_tree_add_14_36_groupi_g52432 (.a(csa_tree_add_14_36_groupi_n_567), .b(csa_tree_add_14_36_groupi_n_381), .y(csa_tree_add_14_36_groupi_n_732));
nand2 csa_tree_add_14_36_groupi_g52433 (.a(csa_tree_add_14_36_groupi_n_568), .b(csa_tree_add_14_36_groupi_n_341), .y(csa_tree_add_14_36_groupi_n_731));
nand2 csa_tree_add_14_36_groupi_g52434 (.a(csa_tree_add_14_36_groupi_n_515), .b(csa_tree_add_14_36_groupi_n_349), .y(csa_tree_add_14_36_groupi_n_730));
nand2 csa_tree_add_14_36_groupi_g52435 (.a(csa_tree_add_14_36_groupi_n_642), .b(csa_tree_add_14_36_groupi_n_325), .y(csa_tree_add_14_36_groupi_n_729));
xor2 csa_tree_add_14_36_groupi_g52436 (.a(n_85), .b(csa_tree_add_14_36_groupi_n_2036), .y(csa_tree_add_14_36_groupi_n_728));
nor2 csa_tree_add_14_36_groupi_g52437 (.a(csa_tree_add_14_36_groupi_n_575), .b(csa_tree_add_14_36_groupi_n_320), .y(csa_tree_add_14_36_groupi_n_727));
nand2 csa_tree_add_14_36_groupi_g52438 (.a(csa_tree_add_14_36_groupi_n_527), .b(csa_tree_add_14_36_groupi_n_344), .y(csa_tree_add_14_36_groupi_n_726));
nand2 csa_tree_add_14_36_groupi_g52439 (.a(csa_tree_add_14_36_groupi_n_523), .b(csa_tree_add_14_36_groupi_n_347), .y(csa_tree_add_14_36_groupi_n_725));
nand2 csa_tree_add_14_36_groupi_g52440 (.a(csa_tree_add_14_36_groupi_n_555), .b(csa_tree_add_14_36_groupi_n_419), .y(csa_tree_add_14_36_groupi_n_724));
nand2 csa_tree_add_14_36_groupi_g52441 (.a(csa_tree_add_14_36_groupi_n_548), .b(csa_tree_add_14_36_groupi_n_346), .y(csa_tree_add_14_36_groupi_n_723));
nand2 csa_tree_add_14_36_groupi_g52442 (.a(csa_tree_add_14_36_groupi_n_519), .b(csa_tree_add_14_36_groupi_n_334), .y(csa_tree_add_14_36_groupi_n_722));
nand2 csa_tree_add_14_36_groupi_g52443 (.a(csa_tree_add_14_36_groupi_n_563), .b(csa_tree_add_14_36_groupi_n_348), .y(csa_tree_add_14_36_groupi_n_721));
nand2 csa_tree_add_14_36_groupi_g52444 (.a(csa_tree_add_14_36_groupi_n_552), .b(csa_tree_add_14_36_groupi_n_387), .y(csa_tree_add_14_36_groupi_n_720));
nand2 csa_tree_add_14_36_groupi_g52445 (.a(csa_tree_add_14_36_groupi_n_545), .b(csa_tree_add_14_36_groupi_n_324), .y(csa_tree_add_14_36_groupi_n_719));
nand2 csa_tree_add_14_36_groupi_g52446 (.a(csa_tree_add_14_36_groupi_n_574), .b(csa_tree_add_14_36_groupi_n_422), .y(csa_tree_add_14_36_groupi_n_718));
nand2 csa_tree_add_14_36_groupi_g52447 (.a(csa_tree_add_14_36_groupi_n_553), .b(csa_tree_add_14_36_groupi_n_377), .y(csa_tree_add_14_36_groupi_n_717));
nand2 csa_tree_add_14_36_groupi_g52448 (.a(csa_tree_add_14_36_groupi_n_641), .b(csa_tree_add_14_36_groupi_n_378), .y(csa_tree_add_14_36_groupi_n_716));
nand2 csa_tree_add_14_36_groupi_g52449 (.a(csa_tree_add_14_36_groupi_n_578), .b(csa_tree_add_14_36_groupi_n_373), .y(csa_tree_add_14_36_groupi_n_715));
nand2 csa_tree_add_14_36_groupi_g52450 (.a(csa_tree_add_14_36_groupi_n_556), .b(csa_tree_add_14_36_groupi_n_391), .y(csa_tree_add_14_36_groupi_n_714));
nand2 csa_tree_add_14_36_groupi_g52451 (.a(csa_tree_add_14_36_groupi_n_571), .b(csa_tree_add_14_36_groupi_n_416), .y(csa_tree_add_14_36_groupi_n_713));
nand2 csa_tree_add_14_36_groupi_g52452 (.a(csa_tree_add_14_36_groupi_n_549), .b(csa_tree_add_14_36_groupi_n_386), .y(csa_tree_add_14_36_groupi_n_712));
nand2 csa_tree_add_14_36_groupi_g52453 (.a(csa_tree_add_14_36_groupi_n_530), .b(csa_tree_add_14_36_groupi_n_317), .y(csa_tree_add_14_36_groupi_n_711));
nand2 csa_tree_add_14_36_groupi_g52454 (.a(csa_tree_add_14_36_groupi_n_566), .b(csa_tree_add_14_36_groupi_n_383), .y(csa_tree_add_14_36_groupi_n_709));
nand2 csa_tree_add_14_36_groupi_g52455 (.a(csa_tree_add_14_36_groupi_n_557), .b(csa_tree_add_14_36_groupi_n_390), .y(csa_tree_add_14_36_groupi_n_708));
nand2 csa_tree_add_14_36_groupi_g52456 (.a(csa_tree_add_14_36_groupi_n_561), .b(csa_tree_add_14_36_groupi_n_388), .y(csa_tree_add_14_36_groupi_n_707));
nand2 csa_tree_add_14_36_groupi_g52457 (.a(csa_tree_add_14_36_groupi_n_562), .b(csa_tree_add_14_36_groupi_n_484), .y(csa_tree_add_14_36_groupi_n_706));
nand2 csa_tree_add_14_36_groupi_g52458 (.a(csa_tree_add_14_36_groupi_n_576), .b(csa_tree_add_14_36_groupi_n_415), .y(csa_tree_add_14_36_groupi_n_705));
nand2 csa_tree_add_14_36_groupi_g52459 (.a(csa_tree_add_14_36_groupi_n_546), .b(csa_tree_add_14_36_groupi_n_382), .y(csa_tree_add_14_36_groupi_n_704));
nand2 csa_tree_add_14_36_groupi_g52460 (.a(csa_tree_add_14_36_groupi_n_573), .b(csa_tree_add_14_36_groupi_n_417), .y(csa_tree_add_14_36_groupi_n_703));
nand2 csa_tree_add_14_36_groupi_g52461 (.a(csa_tree_add_14_36_groupi_n_564), .b(csa_tree_add_14_36_groupi_n_420), .y(csa_tree_add_14_36_groupi_n_702));
inv csa_tree_add_14_36_groupi_g52462 (.a(csa_tree_add_14_36_groupi_n_613), .y(csa_tree_add_14_36_groupi_n_662));
inv csa_tree_add_14_36_groupi_g52463 (.a(csa_tree_add_14_36_groupi_n_2026), .y(csa_tree_add_14_36_groupi_n_661));
inv csa_tree_add_14_36_groupi_g52464 (.a(csa_tree_add_14_36_groupi_n_2051), .y(csa_tree_add_14_36_groupi_n_660));
inv csa_tree_add_14_36_groupi_g52465 (.a(csa_tree_add_14_36_groupi_n_2153), .y(csa_tree_add_14_36_groupi_n_658));
inv csa_tree_add_14_36_groupi_g52466 (.a(csa_tree_add_14_36_groupi_n_2156), .y(csa_tree_add_14_36_groupi_n_657));
inv csa_tree_add_14_36_groupi_g52467 (.a(csa_tree_add_14_36_groupi_n_2124), .y(csa_tree_add_14_36_groupi_n_656));
inv csa_tree_add_14_36_groupi_g52468 (.a(csa_tree_add_14_36_groupi_n_2260), .y(csa_tree_add_14_36_groupi_n_655));
inv csa_tree_add_14_36_groupi_g52469 (.a(csa_tree_add_14_36_groupi_n_2157), .y(csa_tree_add_14_36_groupi_n_654));
inv csa_tree_add_14_36_groupi_g52470 (.a(csa_tree_add_14_36_groupi_n_2154), .y(csa_tree_add_14_36_groupi_n_653));
nand2 csa_tree_add_14_36_groupi_g52472 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_162), .y(csa_tree_add_14_36_groupi_n_649));
nand2 csa_tree_add_14_36_groupi_g52473 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_205), .y(csa_tree_add_14_36_groupi_n_648));
nand2 csa_tree_add_14_36_groupi_g52474 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_311), .y(csa_tree_add_14_36_groupi_n_647));
nand2 csa_tree_add_14_36_groupi_g52475 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_213), .y(csa_tree_add_14_36_groupi_n_646));
nand2 csa_tree_add_14_36_groupi_g52476 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_220), .y(csa_tree_add_14_36_groupi_n_645));
nand2 csa_tree_add_14_36_groupi_g52477 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_226), .y(csa_tree_add_14_36_groupi_n_644));
nand2 csa_tree_add_14_36_groupi_g52478 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_189), .y(csa_tree_add_14_36_groupi_n_643));
nand2 csa_tree_add_14_36_groupi_g52479 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_190), .y(csa_tree_add_14_36_groupi_n_642));
nand2 csa_tree_add_14_36_groupi_g52480 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_299), .y(csa_tree_add_14_36_groupi_n_641));
nand2 csa_tree_add_14_36_groupi_g52481 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_282), .y(csa_tree_add_14_36_groupi_n_640));
nand2 csa_tree_add_14_36_groupi_g52482 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_201), .y(csa_tree_add_14_36_groupi_n_639));
nand2 csa_tree_add_14_36_groupi_g52483 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_195), .y(csa_tree_add_14_36_groupi_n_638));
nor2 csa_tree_add_14_36_groupi_g52484 (.a(csa_tree_add_14_36_groupi_n_492), .b(csa_tree_add_14_36_groupi_n_249), .y(csa_tree_add_14_36_groupi_n_637));
nand2 csa_tree_add_14_36_groupi_g52485 (.a(csa_tree_add_14_36_groupi_n_486), .b(csa_tree_add_14_36_groupi_n_127), .y(csa_tree_add_14_36_groupi_n_636));
nor2 csa_tree_add_14_36_groupi_g52486 (.a(n_2576), .b(csa_tree_add_14_36_groupi_n_251), .y(csa_tree_add_14_36_groupi_n_635));
nand2 csa_tree_add_14_36_groupi_g52487 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_286), .y(csa_tree_add_14_36_groupi_n_634));
nand2 csa_tree_add_14_36_groupi_g52488 (.a(csa_tree_add_14_36_groupi_n_368), .b(csa_tree_add_14_36_groupi_n_481), .y(csa_tree_add_14_36_groupi_n_633));
nand2 csa_tree_add_14_36_groupi_g52489 (.a(csa_tree_add_14_36_groupi_n_359), .b(csa_tree_add_14_36_groupi_n_478), .y(csa_tree_add_14_36_groupi_n_632));
nand2 csa_tree_add_14_36_groupi_g52490 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_152), .y(csa_tree_add_14_36_groupi_n_631));
nand2 csa_tree_add_14_36_groupi_g52491 (.a(csa_tree_add_14_36_groupi_n_364), .b(csa_tree_add_14_36_groupi_n_479), .y(csa_tree_add_14_36_groupi_n_630));
nand2 csa_tree_add_14_36_groupi_g52492 (.a(csa_tree_add_14_36_groupi_n_358), .b(csa_tree_add_14_36_groupi_n_480), .y(csa_tree_add_14_36_groupi_n_629));
nand2 csa_tree_add_14_36_groupi_g52493 (.a(csa_tree_add_14_36_groupi_n_363), .b(csa_tree_add_14_36_groupi_n_475), .y(csa_tree_add_14_36_groupi_n_628));
nand2 csa_tree_add_14_36_groupi_g52494 (.a(csa_tree_add_14_36_groupi_n_365), .b(csa_tree_add_14_36_groupi_n_473), .y(csa_tree_add_14_36_groupi_n_627));
nand2 csa_tree_add_14_36_groupi_g52495 (.a(csa_tree_add_14_36_groupi_n_362), .b(csa_tree_add_14_36_groupi_n_472), .y(csa_tree_add_14_36_groupi_n_626));
nand2 csa_tree_add_14_36_groupi_g52496 (.a(csa_tree_add_14_36_groupi_n_361), .b(csa_tree_add_14_36_groupi_n_471), .y(csa_tree_add_14_36_groupi_n_625));
nand2 csa_tree_add_14_36_groupi_g52497 (.a(csa_tree_add_14_36_groupi_n_370), .b(csa_tree_add_14_36_groupi_n_476), .y(csa_tree_add_14_36_groupi_n_624));
nand2 csa_tree_add_14_36_groupi_g52498 (.a(csa_tree_add_14_36_groupi_n_371), .b(csa_tree_add_14_36_groupi_n_474), .y(csa_tree_add_14_36_groupi_n_623));
nand2 csa_tree_add_14_36_groupi_g52499 (.a(csa_tree_add_14_36_groupi_n_360), .b(csa_tree_add_14_36_groupi_n_468), .y(csa_tree_add_14_36_groupi_n_622));
nand2 csa_tree_add_14_36_groupi_g52500 (.a(csa_tree_add_14_36_groupi_n_369), .b(csa_tree_add_14_36_groupi_n_469), .y(csa_tree_add_14_36_groupi_n_621));
nand2 csa_tree_add_14_36_groupi_g52501 (.a(csa_tree_add_14_36_groupi_n_372), .b(csa_tree_add_14_36_groupi_n_467), .y(csa_tree_add_14_36_groupi_n_620));
nand2 csa_tree_add_14_36_groupi_g52502 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_171), .y(csa_tree_add_14_36_groupi_n_619));
nand2 csa_tree_add_14_36_groupi_g52503 (.a(csa_tree_add_14_36_groupi_n_409), .b(n_2526), .y(csa_tree_add_14_36_groupi_n_618));
nand2 csa_tree_add_14_36_groupi_g52504 (.a(csa_tree_add_14_36_groupi_n_487), .b(n_145), .y(csa_tree_add_14_36_groupi_n_617));
nand2 csa_tree_add_14_36_groupi_g52506 (.a(csa_tree_add_14_36_groupi_n_237), .b(csa_tree_add_14_36_groupi_n_470), .y(csa_tree_add_14_36_groupi_n_615));
nand2 csa_tree_add_14_36_groupi_g52507 (.a(csa_tree_add_14_36_groupi_n_466), .b(csa_tree_add_14_36_groupi_n_255), .y(csa_tree_add_14_36_groupi_n_614));
nor2 csa_tree_add_14_36_groupi_g52508 (.a(csa_tree_add_14_36_groupi_n_408), .b(a_1), .y(csa_tree_add_14_36_groupi_n_613));
nand2 csa_tree_add_14_36_groupi_g52509 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_173), .y(csa_tree_add_14_36_groupi_n_612));
nand2 csa_tree_add_14_36_groupi_g52510 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_174), .y(csa_tree_add_14_36_groupi_n_611));
nand2 csa_tree_add_14_36_groupi_g52511 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_172), .y(csa_tree_add_14_36_groupi_n_610));
nand2 csa_tree_add_14_36_groupi_g52512 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_180), .y(csa_tree_add_14_36_groupi_n_609));
nand2 csa_tree_add_14_36_groupi_g52513 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_179), .y(csa_tree_add_14_36_groupi_n_608));
nand2 csa_tree_add_14_36_groupi_g52514 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_169), .y(csa_tree_add_14_36_groupi_n_607));
nand2 csa_tree_add_14_36_groupi_g52515 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_182), .y(csa_tree_add_14_36_groupi_n_606));
nand2 csa_tree_add_14_36_groupi_g52516 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_158), .y(csa_tree_add_14_36_groupi_n_605));
nand2 csa_tree_add_14_36_groupi_g52517 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_177), .y(csa_tree_add_14_36_groupi_n_604));
nand2 csa_tree_add_14_36_groupi_g52518 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_175), .y(csa_tree_add_14_36_groupi_n_603));
nand2 csa_tree_add_14_36_groupi_g52519 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_157), .y(csa_tree_add_14_36_groupi_n_602));
nand2 csa_tree_add_14_36_groupi_g52520 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_168), .y(csa_tree_add_14_36_groupi_n_601));
nand2 csa_tree_add_14_36_groupi_g52521 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_156), .y(csa_tree_add_14_36_groupi_n_600));
nand2 csa_tree_add_14_36_groupi_g52522 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_155), .y(csa_tree_add_14_36_groupi_n_599));
nand2 csa_tree_add_14_36_groupi_g52523 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_159), .y(csa_tree_add_14_36_groupi_n_598));
nand2 csa_tree_add_14_36_groupi_g52524 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_166), .y(csa_tree_add_14_36_groupi_n_597));
nand2 csa_tree_add_14_36_groupi_g52525 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_165), .y(csa_tree_add_14_36_groupi_n_596));
nand2 csa_tree_add_14_36_groupi_g52526 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_181), .y(csa_tree_add_14_36_groupi_n_595));
nand2 csa_tree_add_14_36_groupi_g52527 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_139), .y(csa_tree_add_14_36_groupi_n_594));
nand2 csa_tree_add_14_36_groupi_g52528 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_154), .y(csa_tree_add_14_36_groupi_n_593));
nand2 csa_tree_add_14_36_groupi_g52529 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_161), .y(csa_tree_add_14_36_groupi_n_592));
nand2 csa_tree_add_14_36_groupi_g52530 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_176), .y(csa_tree_add_14_36_groupi_n_591));
nand2 csa_tree_add_14_36_groupi_g52531 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_164), .y(csa_tree_add_14_36_groupi_n_590));
nand2 csa_tree_add_14_36_groupi_g52532 (.a(csa_tree_add_14_36_groupi_n_399), .b(csa_tree_add_14_36_groupi_n_167), .y(csa_tree_add_14_36_groupi_n_589));
nand2 csa_tree_add_14_36_groupi_g52533 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_160), .y(csa_tree_add_14_36_groupi_n_588));
nand2 csa_tree_add_14_36_groupi_g52534 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_153), .y(csa_tree_add_14_36_groupi_n_587));
nand2 csa_tree_add_14_36_groupi_g52535 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_142), .y(csa_tree_add_14_36_groupi_n_586));
nand2 csa_tree_add_14_36_groupi_g52536 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_178), .y(csa_tree_add_14_36_groupi_n_585));
nand2 csa_tree_add_14_36_groupi_g52537 (.a(csa_tree_add_14_36_groupi_n_403), .b(csa_tree_add_14_36_groupi_n_151), .y(csa_tree_add_14_36_groupi_n_584));
nand2 csa_tree_add_14_36_groupi_g52551 (.a(csa_tree_add_14_36_groupi_n_367), .b(csa_tree_add_14_36_groupi_n_95), .y(csa_tree_add_14_36_groupi_n_651));
nand2 csa_tree_add_14_36_groupi_g52552 (.a(csa_tree_add_14_36_groupi_n_366), .b(csa_tree_add_14_36_groupi_n_477), .y(csa_tree_add_14_36_groupi_n_650));
inv csa_tree_add_14_36_groupi_g52553 (.a(csa_tree_add_14_36_groupi_n_582), .y(csa_tree_add_14_36_groupi_n_583));
nand2 csa_tree_add_14_36_groupi_g52554 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_199), .y(csa_tree_add_14_36_groupi_n_581));
nand2 csa_tree_add_14_36_groupi_g52555 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_141), .y(csa_tree_add_14_36_groupi_n_580));
nand2 csa_tree_add_14_36_groupi_g52556 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_252), .y(csa_tree_add_14_36_groupi_n_579));
nand2 csa_tree_add_14_36_groupi_g52557 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_221), .y(csa_tree_add_14_36_groupi_n_578));
nand2 csa_tree_add_14_36_groupi_g52558 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_294), .y(csa_tree_add_14_36_groupi_n_577));
nand2 csa_tree_add_14_36_groupi_g52559 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_276), .y(csa_tree_add_14_36_groupi_n_576));
nor2 csa_tree_add_14_36_groupi_g52560 (.a(csa_tree_add_14_36_groupi_n_406), .b(csa_tree_add_14_36_groupi_n_163), .y(csa_tree_add_14_36_groupi_n_575));
nand2 csa_tree_add_14_36_groupi_g52561 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_218), .y(csa_tree_add_14_36_groupi_n_574));
nand2 csa_tree_add_14_36_groupi_g52562 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_266), .y(csa_tree_add_14_36_groupi_n_573));
nand2 csa_tree_add_14_36_groupi_g52563 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_267), .y(csa_tree_add_14_36_groupi_n_572));
nand2 csa_tree_add_14_36_groupi_g52564 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_296), .y(csa_tree_add_14_36_groupi_n_571));
nand2 csa_tree_add_14_36_groupi_g52565 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_281), .y(csa_tree_add_14_36_groupi_n_570));
nand2 csa_tree_add_14_36_groupi_g52566 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_207), .y(csa_tree_add_14_36_groupi_n_569));
nand2 csa_tree_add_14_36_groupi_g52567 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_271), .y(csa_tree_add_14_36_groupi_n_568));
nand2 csa_tree_add_14_36_groupi_g52568 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_200), .y(csa_tree_add_14_36_groupi_n_567));
nand2 csa_tree_add_14_36_groupi_g52569 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_202), .y(csa_tree_add_14_36_groupi_n_566));
nand2 csa_tree_add_14_36_groupi_g52570 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_280), .y(csa_tree_add_14_36_groupi_n_565));
nand2 csa_tree_add_14_36_groupi_g52571 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_209), .y(csa_tree_add_14_36_groupi_n_564));
nand2 csa_tree_add_14_36_groupi_g52572 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_268), .y(csa_tree_add_14_36_groupi_n_563));
nand2 csa_tree_add_14_36_groupi_g52573 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_309), .y(csa_tree_add_14_36_groupi_n_562));
nand2 csa_tree_add_14_36_groupi_g52574 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_208), .y(csa_tree_add_14_36_groupi_n_561));
nand2 csa_tree_add_14_36_groupi_g52575 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_194), .y(csa_tree_add_14_36_groupi_n_560));
nand2 csa_tree_add_14_36_groupi_g52576 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_140), .y(csa_tree_add_14_36_groupi_n_559));
nand2 csa_tree_add_14_36_groupi_g52577 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_265), .y(csa_tree_add_14_36_groupi_n_558));
nand2 csa_tree_add_14_36_groupi_g52578 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_206), .y(csa_tree_add_14_36_groupi_n_557));
nand2 csa_tree_add_14_36_groupi_g52579 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_197), .y(csa_tree_add_14_36_groupi_n_556));
nand2 csa_tree_add_14_36_groupi_g52580 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_193), .y(csa_tree_add_14_36_groupi_n_555));
nand2 csa_tree_add_14_36_groupi_g52581 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_216), .y(csa_tree_add_14_36_groupi_n_554));
nand2 csa_tree_add_14_36_groupi_g52582 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_312), .y(csa_tree_add_14_36_groupi_n_553));
nand2 csa_tree_add_14_36_groupi_g52583 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_273), .y(csa_tree_add_14_36_groupi_n_552));
nand2 csa_tree_add_14_36_groupi_g52584 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_191), .y(csa_tree_add_14_36_groupi_n_551));
nand2 csa_tree_add_14_36_groupi_g52585 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_297), .y(csa_tree_add_14_36_groupi_n_550));
nand2 csa_tree_add_14_36_groupi_g52586 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_214), .y(csa_tree_add_14_36_groupi_n_549));
nand2 csa_tree_add_14_36_groupi_g52587 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_184), .y(csa_tree_add_14_36_groupi_n_548));
nand2 csa_tree_add_14_36_groupi_g52588 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_275), .y(csa_tree_add_14_36_groupi_n_547));
nand2 csa_tree_add_14_36_groupi_g52589 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_224), .y(csa_tree_add_14_36_groupi_n_546));
nand2 csa_tree_add_14_36_groupi_g52590 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_192), .y(csa_tree_add_14_36_groupi_n_545));
nand2 csa_tree_add_14_36_groupi_g52591 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_198), .y(csa_tree_add_14_36_groupi_n_544));
nand2 csa_tree_add_14_36_groupi_g52592 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_225), .y(csa_tree_add_14_36_groupi_n_543));
nand2 csa_tree_add_14_36_groupi_g52593 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_284), .y(csa_tree_add_14_36_groupi_n_542));
nand2 csa_tree_add_14_36_groupi_g52594 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_212), .y(csa_tree_add_14_36_groupi_n_541));
nand2 csa_tree_add_14_36_groupi_g52595 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_285), .y(csa_tree_add_14_36_groupi_n_540));
nand2 csa_tree_add_14_36_groupi_g52596 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_272), .y(csa_tree_add_14_36_groupi_n_539));
nand2 csa_tree_add_14_36_groupi_g52597 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_279), .y(csa_tree_add_14_36_groupi_n_538));
nand2 csa_tree_add_14_36_groupi_g52598 (.a(csa_tree_add_14_36_groupi_n_397), .b(csa_tree_add_14_36_groupi_n_217), .y(csa_tree_add_14_36_groupi_n_537));
nand2 csa_tree_add_14_36_groupi_g52599 (.a(csa_tree_add_14_36_groupi_n_395), .b(csa_tree_add_14_36_groupi_n_196), .y(csa_tree_add_14_36_groupi_n_536));
nand2 csa_tree_add_14_36_groupi_g52600 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_223), .y(csa_tree_add_14_36_groupi_n_535));
nand2 csa_tree_add_14_36_groupi_g52601 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_277), .y(csa_tree_add_14_36_groupi_n_534));
nand2 csa_tree_add_14_36_groupi_g52602 (.a(csa_tree_add_14_36_groupi_n_401), .b(csa_tree_add_14_36_groupi_n_187), .y(csa_tree_add_14_36_groupi_n_533));
nand2 csa_tree_add_14_36_groupi_g52603 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_288), .y(csa_tree_add_14_36_groupi_n_532));
nand2 csa_tree_add_14_36_groupi_g52604 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_287), .y(csa_tree_add_14_36_groupi_n_531));
nand2 csa_tree_add_14_36_groupi_g52605 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_290), .y(csa_tree_add_14_36_groupi_n_530));
nand2 csa_tree_add_14_36_groupi_g52606 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_289), .y(csa_tree_add_14_36_groupi_n_529));
nor2 csa_tree_add_14_36_groupi_g52607 (.a(csa_tree_add_14_36_groupi_n_483), .b(csa_tree_add_14_36_groupi_n_75), .y(csa_tree_add_14_36_groupi_n_528));
nand2 csa_tree_add_14_36_groupi_g52608 (.a(csa_tree_add_14_36_groupi_n_407), .b(csa_tree_add_14_36_groupi_n_234), .y(csa_tree_add_14_36_groupi_n_527));
nor2 csa_tree_add_14_36_groupi_g52609 (.a(csa_tree_add_14_36_groupi_n_482), .b(csa_tree_add_14_36_groupi_n_59), .y(csa_tree_add_14_36_groupi_n_526));
nand2 csa_tree_add_14_36_groupi_g52610 (.a(csa_tree_add_14_36_groupi_n_404), .b(b_15), .y(csa_tree_add_14_36_groupi_n_525));
nand2 csa_tree_add_14_36_groupi_g52611 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_306), .y(csa_tree_add_14_36_groupi_n_524));
nand2 csa_tree_add_14_36_groupi_g52612 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_302), .y(csa_tree_add_14_36_groupi_n_523));
nand2 csa_tree_add_14_36_groupi_g52613 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_301), .y(csa_tree_add_14_36_groupi_n_522));
nand2 csa_tree_add_14_36_groupi_g52614 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_305), .y(csa_tree_add_14_36_groupi_n_521));
nand2 csa_tree_add_14_36_groupi_g52615 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_303), .y(csa_tree_add_14_36_groupi_n_520));
nand2 csa_tree_add_14_36_groupi_g52616 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_308), .y(csa_tree_add_14_36_groupi_n_519));
nor2 csa_tree_add_14_36_groupi_g52617 (.a(csa_tree_add_14_36_groupi_n_405), .b(csa_tree_add_14_36_groupi_n_235), .y(csa_tree_add_14_36_groupi_n_518));
nand2 csa_tree_add_14_36_groupi_g52618 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_307), .y(csa_tree_add_14_36_groupi_n_517));
nand2 csa_tree_add_14_36_groupi_g52619 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_304), .y(csa_tree_add_14_36_groupi_n_516));
nand2 csa_tree_add_14_36_groupi_g52620 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_300), .y(csa_tree_add_14_36_groupi_n_515));
nand2 csa_tree_add_14_36_groupi_g52622 (.a(csa_tree_add_14_36_groupi_n_404), .b(csa_tree_add_14_36_groupi_n_310), .y(csa_tree_add_14_36_groupi_n_513));
xor2 csa_tree_add_14_36_groupi_g52628 (.a(n_86), .b(csa_tree_add_14_36_groupi_n_2066), .y(result_0__0_));
xor2 csa_tree_add_14_36_groupi_g52629 (.a(n_123), .b(csa_tree_add_14_36_groupi_n_2027), .y(csa_tree_add_14_36_groupi_n_507));
xor2 csa_tree_add_14_36_groupi_g52630 (.a(n_139), .b(csa_tree_add_14_36_groupi_n_2155), .y(csa_tree_add_14_36_groupi_n_506));
xor2 csa_tree_add_14_36_groupi_g52631 (.a(n_145), .b(csa_tree_add_14_36_groupi_n_2158), .y(csa_tree_add_14_36_groupi_n_505));
xor2 csa_tree_add_14_36_groupi_g52632 (.a(n_127), .b(csa_tree_add_14_36_groupi_n_2034), .y(csa_tree_add_14_36_groupi_n_504));
xor2 csa_tree_add_14_36_groupi_g52633 (.a(csa_tree_add_14_36_groupi_n_136), .b(csa_tree_add_14_36_groupi_n_2028), .y(csa_tree_add_14_36_groupi_n_582));
xor2 csa_tree_add_14_36_groupi_g52634 (.a(n_135), .b(csa_tree_add_14_36_groupi_n_2304), .y(csa_tree_add_14_36_groupi_n_503));
xor2 csa_tree_add_14_36_groupi_g52635 (.a(n_149), .b(csa_tree_add_14_36_groupi_n_2035), .y(csa_tree_add_14_36_groupi_n_502));
inv csa_tree_add_14_36_groupi_g52636 (.a(csa_tree_add_14_36_groupi_n_491), .y(csa_tree_add_14_36_groupi_n_501));
inv csa_tree_add_14_36_groupi_g52637 (.a(csa_tree_add_14_36_groupi_n_489), .y(csa_tree_add_14_36_groupi_n_500));
inv csa_tree_add_14_36_groupi_g52638 (.a(csa_tree_add_14_36_groupi_n_454), .y(csa_tree_add_14_36_groupi_n_499));
inv csa_tree_add_14_36_groupi_g52639 (.a(csa_tree_add_14_36_groupi_n_497), .y(csa_tree_add_14_36_groupi_n_498));
nand2 csa_tree_add_14_36_groupi_g52640 (.a(csa_tree_add_14_36_groupi_n_151), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_496));
nand2 csa_tree_add_14_36_groupi_g52641 (.a(csa_tree_add_14_36_groupi_n_250), .b(csa_tree_add_14_36_groupi_n_292), .y(csa_tree_add_14_36_groupi_n_495));
nand2 csa_tree_add_14_36_groupi_g52643 (.a(csa_tree_add_14_36_groupi_n_217), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_493));
nor2 csa_tree_add_14_36_groupi_g52644 (.a(csa_tree_add_14_36_groupi_n_292), .b(a_1), .y(csa_tree_add_14_36_groupi_n_492));
nor2 csa_tree_add_14_36_groupi_g52645 (.a(csa_tree_add_14_36_groupi_n_247), .b(csa_tree_add_14_36_groupi_n_253), .y(csa_tree_add_14_36_groupi_n_491));
nand2 csa_tree_add_14_36_groupi_g52646 (.a(csa_tree_add_14_36_groupi_n_248), .b(n_2577), .y(csa_tree_add_14_36_groupi_n_490));
nor2 csa_tree_add_14_36_groupi_g52647 (.a(csa_tree_add_14_36_groupi_n_245), .b(csa_tree_add_14_36_groupi_n_242), .y(csa_tree_add_14_36_groupi_n_489));
nand2 csa_tree_add_14_36_groupi_g52648 (.a(csa_tree_add_14_36_groupi_n_197), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_488));
nand2 csa_tree_add_14_36_groupi_g52649 (.a(csa_tree_add_14_36_groupi_n_63), .b(csa_tree_add_14_36_groupi_n_2028), .y(csa_tree_add_14_36_groupi_n_487));
nor2 csa_tree_add_14_36_groupi_g52650 (.a(csa_tree_add_14_36_groupi_n_129), .b(csa_tree_add_14_36_groupi_n_269), .y(csa_tree_add_14_36_groupi_n_486));
nand2 csa_tree_add_14_36_groupi_g52651 (.a(n_137), .b(csa_tree_add_14_36_groupi_n_264), .y(csa_tree_add_14_36_groupi_n_485));
nand2 csa_tree_add_14_36_groupi_g52652 (.a(csa_tree_add_14_36_groupi_n_192), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_484));
nor2 csa_tree_add_14_36_groupi_g52653 (.a(n_2451), .b(csa_tree_add_14_36_groupi_n_121), .y(csa_tree_add_14_36_groupi_n_483));
nor2 csa_tree_add_14_36_groupi_g52654 (.a(csa_tree_add_14_36_groupi_n_241), .b(csa_tree_add_14_36_groupi_n_117), .y(csa_tree_add_14_36_groupi_n_482));
nand2 csa_tree_add_14_36_groupi_g52655 (.a(csa_tree_add_14_36_groupi_n_183), .b(b_0), .y(csa_tree_add_14_36_groupi_n_481));
nand2 csa_tree_add_14_36_groupi_g52656 (.a(csa_tree_add_14_36_groupi_n_186), .b(b_0), .y(csa_tree_add_14_36_groupi_n_480));
nand2 csa_tree_add_14_36_groupi_g52657 (.a(csa_tree_add_14_36_groupi_n_215), .b(b_0), .y(csa_tree_add_14_36_groupi_n_479));
nand2 csa_tree_add_14_36_groupi_g52658 (.a(csa_tree_add_14_36_groupi_n_211), .b(b_0), .y(csa_tree_add_14_36_groupi_n_478));
nand2 csa_tree_add_14_36_groupi_g52659 (.a(csa_tree_add_14_36_groupi_n_188), .b(b_0), .y(csa_tree_add_14_36_groupi_n_477));
nand2 csa_tree_add_14_36_groupi_g52660 (.a(csa_tree_add_14_36_groupi_n_222), .b(b_0), .y(csa_tree_add_14_36_groupi_n_476));
nand2 csa_tree_add_14_36_groupi_g52661 (.a(csa_tree_add_14_36_groupi_n_283), .b(b_0), .y(csa_tree_add_14_36_groupi_n_475));
nand2 csa_tree_add_14_36_groupi_g52662 (.a(csa_tree_add_14_36_groupi_n_274), .b(b_0), .y(csa_tree_add_14_36_groupi_n_474));
nand2 csa_tree_add_14_36_groupi_g52663 (.a(csa_tree_add_14_36_groupi_n_185), .b(b_0), .y(csa_tree_add_14_36_groupi_n_473));
nand2 csa_tree_add_14_36_groupi_g52664 (.a(csa_tree_add_14_36_groupi_n_219), .b(b_0), .y(csa_tree_add_14_36_groupi_n_472));
nand2 csa_tree_add_14_36_groupi_g52665 (.a(csa_tree_add_14_36_groupi_n_278), .b(b_0), .y(csa_tree_add_14_36_groupi_n_471));
nand2 csa_tree_add_14_36_groupi_g52666 (.a(csa_tree_add_14_36_groupi_n_203), .b(b_0), .y(csa_tree_add_14_36_groupi_n_470));
nand2 csa_tree_add_14_36_groupi_g52667 (.a(csa_tree_add_14_36_groupi_n_170), .b(b_0), .y(csa_tree_add_14_36_groupi_n_469));
nand2 csa_tree_add_14_36_groupi_g52668 (.a(csa_tree_add_14_36_groupi_n_270), .b(b_0), .y(csa_tree_add_14_36_groupi_n_468));
nand2 csa_tree_add_14_36_groupi_g52669 (.a(csa_tree_add_14_36_groupi_n_210), .b(b_0), .y(csa_tree_add_14_36_groupi_n_467));
nor2 csa_tree_add_14_36_groupi_g52670 (.a(csa_tree_add_14_36_groupi_n_204), .b(csa_tree_add_14_36_groupi_n_293), .y(csa_tree_add_14_36_groupi_n_466));
nor2 csa_tree_add_14_36_groupi_g52671 (.a(csa_tree_add_14_36_groupi_n_134), .b(csa_tree_add_14_36_groupi_n_291), .y(csa_tree_add_14_36_groupi_n_465));
nand2 csa_tree_add_14_36_groupi_g52672 (.a(csa_tree_add_14_36_groupi_n_176), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_464));
nand2 csa_tree_add_14_36_groupi_g52673 (.a(csa_tree_add_14_36_groupi_n_174), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_463));
nand2 csa_tree_add_14_36_groupi_g52674 (.a(csa_tree_add_14_36_groupi_n_180), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_462));
nand2 csa_tree_add_14_36_groupi_g52675 (.a(csa_tree_add_14_36_groupi_n_153), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_461));
nand2 csa_tree_add_14_36_groupi_g52676 (.a(csa_tree_add_14_36_groupi_n_175), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_460));
nand2 csa_tree_add_14_36_groupi_g52677 (.a(csa_tree_add_14_36_groupi_n_173), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_459));
nand2 csa_tree_add_14_36_groupi_g52678 (.a(csa_tree_add_14_36_groupi_n_164), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_458));
nand2 csa_tree_add_14_36_groupi_g52679 (.a(csa_tree_add_14_36_groupi_n_161), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_457));
nand2 csa_tree_add_14_36_groupi_g52680 (.a(csa_tree_add_14_36_groupi_n_157), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_456));
nand2 csa_tree_add_14_36_groupi_g52681 (.a(csa_tree_add_14_36_groupi_n_158), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_455));
nor2 csa_tree_add_14_36_groupi_g52682 (.a(csa_tree_add_14_36_groupi_n_246), .b(csa_tree_add_14_36_groupi_n_243), .y(csa_tree_add_14_36_groupi_n_454));
nand2 csa_tree_add_14_36_groupi_g52683 (.a(csa_tree_add_14_36_groupi_n_165), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_453));
nand2 csa_tree_add_14_36_groupi_g52684 (.a(csa_tree_add_14_36_groupi_n_182), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_452));
nand2 csa_tree_add_14_36_groupi_g52685 (.a(csa_tree_add_14_36_groupi_n_156), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_451));
nand2 csa_tree_add_14_36_groupi_g52686 (.a(csa_tree_add_14_36_groupi_n_169), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_450));
nand2 csa_tree_add_14_36_groupi_g52687 (.a(csa_tree_add_14_36_groupi_n_167), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_449));
nand2 csa_tree_add_14_36_groupi_g52688 (.a(csa_tree_add_14_36_groupi_n_178), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_448));
nand2 csa_tree_add_14_36_groupi_g52689 (.a(csa_tree_add_14_36_groupi_n_166), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_447));
nand2 csa_tree_add_14_36_groupi_g52690 (.a(csa_tree_add_14_36_groupi_n_177), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_446));
nand2 csa_tree_add_14_36_groupi_g52691 (.a(csa_tree_add_14_36_groupi_n_172), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_445));
nand2 csa_tree_add_14_36_groupi_g52692 (.a(csa_tree_add_14_36_groupi_n_155), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_444));
nand2 csa_tree_add_14_36_groupi_g52693 (.a(csa_tree_add_14_36_groupi_n_171), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_443));
nand2 csa_tree_add_14_36_groupi_g52694 (.a(csa_tree_add_14_36_groupi_n_168), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_442));
nand2 csa_tree_add_14_36_groupi_g52695 (.a(csa_tree_add_14_36_groupi_n_159), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_441));
nand2 csa_tree_add_14_36_groupi_g52696 (.a(csa_tree_add_14_36_groupi_n_152), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_440));
nand2 csa_tree_add_14_36_groupi_g52697 (.a(csa_tree_add_14_36_groupi_n_160), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_439));
nand2 csa_tree_add_14_36_groupi_g52698 (.a(csa_tree_add_14_36_groupi_n_154), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_438));
nand2 csa_tree_add_14_36_groupi_g52699 (.a(csa_tree_add_14_36_groupi_n_181), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_437));
nand2 csa_tree_add_14_36_groupi_g52700 (.a(csa_tree_add_14_36_groupi_n_179), .b(csa_tree_add_14_36_groupi_n_144), .y(csa_tree_add_14_36_groupi_n_436));
nand2 csa_tree_add_14_36_groupi_g52701 (.a(csa_tree_add_14_36_groupi_n_162), .b(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_435));
nand2 csa_tree_add_14_36_groupi_g52702 (.a(csa_tree_add_14_36_groupi_n_266), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_434));
nand2 csa_tree_add_14_36_groupi_g52703 (.a(csa_tree_add_14_36_groupi_n_267), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_433));
nand2 csa_tree_add_14_36_groupi_g52704 (.a(csa_tree_add_14_36_groupi_n_280), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_432));
nand2 csa_tree_add_14_36_groupi_g52705 (.a(csa_tree_add_14_36_groupi_n_294), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_431));
nand2 csa_tree_add_14_36_groupi_g52706 (.a(csa_tree_add_14_36_groupi_n_195), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_430));
nand2 csa_tree_add_14_36_groupi_g52707 (.a(csa_tree_add_14_36_groupi_n_194), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_429));
nand2 csa_tree_add_14_36_groupi_g52708 (.a(csa_tree_add_14_36_groupi_n_209), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_428));
nand2 csa_tree_add_14_36_groupi_g52709 (.a(csa_tree_add_14_36_groupi_n_281), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_427));
nand2 csa_tree_add_14_36_groupi_g52710 (.a(csa_tree_add_14_36_groupi_n_198), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_426));
nand2 csa_tree_add_14_36_groupi_g52711 (.a(csa_tree_add_14_36_groupi_n_224), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_425));
nand2 csa_tree_add_14_36_groupi_g52712 (.a(csa_tree_add_14_36_groupi_n_189), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_424));
nand2 csa_tree_add_14_36_groupi_g52713 (.a(csa_tree_add_14_36_groupi_n_311), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_423));
nand2 csa_tree_add_14_36_groupi_g52714 (.a(csa_tree_add_14_36_groupi_n_190), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_422));
nand2 csa_tree_add_14_36_groupi_g52715 (.a(csa_tree_add_14_36_groupi_n_226), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_421));
nand2 csa_tree_add_14_36_groupi_g52716 (.a(csa_tree_add_14_36_groupi_n_214), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_420));
nand2 csa_tree_add_14_36_groupi_g52717 (.a(csa_tree_add_14_36_groupi_n_208), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_419));
nand2 csa_tree_add_14_36_groupi_g52718 (.a(csa_tree_add_14_36_groupi_n_205), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_418));
nand2 csa_tree_add_14_36_groupi_g52719 (.a(csa_tree_add_14_36_groupi_n_200), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_417));
nand2 csa_tree_add_14_36_groupi_g52720 (.a(csa_tree_add_14_36_groupi_n_285), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_416));
nand2 csa_tree_add_14_36_groupi_g52721 (.a(csa_tree_add_14_36_groupi_n_273), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_415));
nand2 csa_tree_add_14_36_groupi_g52722 (.a(csa_tree_add_14_36_groupi_n_225), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_414));
nand2 csa_tree_add_14_36_groupi_g52723 (.a(csa_tree_add_14_36_groupi_n_72), .b(csa_tree_add_14_36_groupi_n_2027), .y(csa_tree_add_14_36_groupi_n_413));
nand2 csa_tree_add_14_36_groupi_g52724 (.a(n_123), .b(csa_tree_add_14_36_groupi_n_295), .y(csa_tree_add_14_36_groupi_n_412));
nand2 csa_tree_add_14_36_groupi_g52726 (.a(n_86), .b(csa_tree_add_14_36_groupi_n_2066), .y(csa_tree_add_14_36_groupi_n_497));
inv csa_tree_add_14_36_groupi_g52727 (.a(csa_tree_add_14_36_groupi_n_351), .y(csa_tree_add_14_36_groupi_n_411));
inv csa_tree_add_14_36_groupi_g52728 (.a(csa_tree_add_14_36_groupi_n_339), .y(csa_tree_add_14_36_groupi_n_410));
inv csa_tree_add_14_36_groupi_g52729 (.a(csa_tree_add_14_36_groupi_n_407), .y(csa_tree_add_14_36_groupi_n_406));
inv csa_tree_add_14_36_groupi_g52730 (.a(csa_tree_add_14_36_groupi_n_404), .y(csa_tree_add_14_36_groupi_n_405));
inv csa_tree_add_14_36_groupi_g52731 (.a(n_2467), .y(csa_tree_add_14_36_groupi_n_403));
inv csa_tree_add_14_36_groupi_g52732 (.a(n_2463), .y(csa_tree_add_14_36_groupi_n_401));
inv csa_tree_add_14_36_groupi_g52733 (.a(n_2678), .y(csa_tree_add_14_36_groupi_n_399));
inv csa_tree_add_14_36_groupi_g52734 (.a(n_2690), .y(csa_tree_add_14_36_groupi_n_397));
inv csa_tree_add_14_36_groupi_g52735 (.a(n_2457), .y(csa_tree_add_14_36_groupi_n_395));
nand2 csa_tree_add_14_36_groupi_g52736 (.a(csa_tree_add_14_36_groupi_n_187), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_393));
nand2 csa_tree_add_14_36_groupi_g52737 (.a(csa_tree_add_14_36_groupi_n_312), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_392));
nand2 csa_tree_add_14_36_groupi_g52738 (.a(csa_tree_add_14_36_groupi_n_193), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_391));
nand2 csa_tree_add_14_36_groupi_g52739 (.a(csa_tree_add_14_36_groupi_n_207), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_390));
nand2 csa_tree_add_14_36_groupi_g52740 (.a(csa_tree_add_14_36_groupi_n_201), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_389));
nand2 csa_tree_add_14_36_groupi_g52741 (.a(csa_tree_add_14_36_groupi_n_212), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_388));
nand2 csa_tree_add_14_36_groupi_g52742 (.a(csa_tree_add_14_36_groupi_n_296), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_387));
nand2 csa_tree_add_14_36_groupi_g52743 (.a(csa_tree_add_14_36_groupi_n_275), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_386));
nand2 csa_tree_add_14_36_groupi_g52744 (.a(csa_tree_add_14_36_groupi_n_279), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_385));
nand2 csa_tree_add_14_36_groupi_g52745 (.a(csa_tree_add_14_36_groupi_n_277), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_384));
nand2 csa_tree_add_14_36_groupi_g52746 (.a(csa_tree_add_14_36_groupi_n_196), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_383));
nand2 csa_tree_add_14_36_groupi_g52747 (.a(csa_tree_add_14_36_groupi_n_221), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_382));
nand2 csa_tree_add_14_36_groupi_g52748 (.a(csa_tree_add_14_36_groupi_n_299), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_381));
nand2 csa_tree_add_14_36_groupi_g52749 (.a(csa_tree_add_14_36_groupi_n_206), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_380));
nand2 csa_tree_add_14_36_groupi_g52750 (.a(csa_tree_add_14_36_groupi_n_272), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_379));
nand2 csa_tree_add_14_36_groupi_g52751 (.a(csa_tree_add_14_36_groupi_n_199), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_378));
nand2 csa_tree_add_14_36_groupi_g52752 (.a(csa_tree_add_14_36_groupi_n_202), .b(csa_tree_add_14_36_groupi_n_257), .y(csa_tree_add_14_36_groupi_n_377));
nand2 csa_tree_add_14_36_groupi_g52753 (.a(csa_tree_add_14_36_groupi_n_218), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_376));
nand2 csa_tree_add_14_36_groupi_g52754 (.a(csa_tree_add_14_36_groupi_n_276), .b(csa_tree_add_14_36_groupi_n_150), .y(csa_tree_add_14_36_groupi_n_375));
nand2 csa_tree_add_14_36_groupi_g52755 (.a(csa_tree_add_14_36_groupi_n_282), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_374));
nand2 csa_tree_add_14_36_groupi_g52756 (.a(csa_tree_add_14_36_groupi_n_309), .b(csa_tree_add_14_36_groupi_n_146), .y(csa_tree_add_14_36_groupi_n_373));
nand2 csa_tree_add_14_36_groupi_g52757 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_222), .y(csa_tree_add_14_36_groupi_n_372));
nand2 csa_tree_add_14_36_groupi_g52758 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_219), .y(csa_tree_add_14_36_groupi_n_371));
nand2 csa_tree_add_14_36_groupi_g52759 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_186), .y(csa_tree_add_14_36_groupi_n_370));
nand2 csa_tree_add_14_36_groupi_g52760 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_183), .y(csa_tree_add_14_36_groupi_n_369));
nand2 csa_tree_add_14_36_groupi_g52761 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_283), .y(csa_tree_add_14_36_groupi_n_368));
nand2 csa_tree_add_14_36_groupi_g52762 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_211), .y(csa_tree_add_14_36_groupi_n_367));
nand2 csa_tree_add_14_36_groupi_g52763 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_170), .y(csa_tree_add_14_36_groupi_n_366));
nand2 csa_tree_add_14_36_groupi_g52764 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_188), .y(csa_tree_add_14_36_groupi_n_365));
nand2 csa_tree_add_14_36_groupi_g52765 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_203), .y(csa_tree_add_14_36_groupi_n_364));
nand2 csa_tree_add_14_36_groupi_g52766 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_210), .y(csa_tree_add_14_36_groupi_n_363));
nand2 csa_tree_add_14_36_groupi_g52767 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_185), .y(csa_tree_add_14_36_groupi_n_362));
nand2 csa_tree_add_14_36_groupi_g52768 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_270), .y(csa_tree_add_14_36_groupi_n_361));
nand2 csa_tree_add_14_36_groupi_g52769 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_274), .y(csa_tree_add_14_36_groupi_n_360));
nand2 csa_tree_add_14_36_groupi_g52770 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_278), .y(csa_tree_add_14_36_groupi_n_359));
nand2 csa_tree_add_14_36_groupi_g52771 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_215), .y(csa_tree_add_14_36_groupi_n_358));
nand2 csa_tree_add_14_36_groupi_g52772 (.a(csa_tree_add_14_36_groupi_n_310), .b(n_2583), .y(csa_tree_add_14_36_groupi_n_357));
nand2 csa_tree_add_14_36_groupi_g52773 (.a(csa_tree_add_14_36_groupi_n_302), .b(n_2583), .y(csa_tree_add_14_36_groupi_n_356));
nand2 csa_tree_add_14_36_groupi_g52774 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_286), .y(csa_tree_add_14_36_groupi_n_355));
nand2 csa_tree_add_14_36_groupi_g52775 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_301), .y(csa_tree_add_14_36_groupi_n_354));
nand2 csa_tree_add_14_36_groupi_g52776 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_297), .y(csa_tree_add_14_36_groupi_n_353));
nand2 csa_tree_add_14_36_groupi_g52777 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_300), .y(csa_tree_add_14_36_groupi_n_352));
nor2 csa_tree_add_14_36_groupi_g52778 (.a(csa_tree_add_14_36_groupi_n_255), .b(csa_tree_add_14_36_groupi_n_163), .y(csa_tree_add_14_36_groupi_n_351));
nand2 csa_tree_add_14_36_groupi_g52779 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_191), .y(csa_tree_add_14_36_groupi_n_350));
nand2 csa_tree_add_14_36_groupi_g52780 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_308), .y(csa_tree_add_14_36_groupi_n_349));
nand2 csa_tree_add_14_36_groupi_g52781 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_213), .y(csa_tree_add_14_36_groupi_n_348));
nand2 csa_tree_add_14_36_groupi_g52782 (.a(csa_tree_add_14_36_groupi_n_303), .b(n_2583), .y(csa_tree_add_14_36_groupi_n_347));
nand2 csa_tree_add_14_36_groupi_g52783 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_284), .y(csa_tree_add_14_36_groupi_n_346));
nand2 csa_tree_add_14_36_groupi_g52784 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_216), .y(csa_tree_add_14_36_groupi_n_345));
nand2 csa_tree_add_14_36_groupi_g52785 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_265), .y(csa_tree_add_14_36_groupi_n_344));
nand2 csa_tree_add_14_36_groupi_g52786 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_184), .y(csa_tree_add_14_36_groupi_n_343));
nand2 csa_tree_add_14_36_groupi_g52787 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_271), .y(csa_tree_add_14_36_groupi_n_342));
nand2 csa_tree_add_14_36_groupi_g52788 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_220), .y(csa_tree_add_14_36_groupi_n_341));
nand2 csa_tree_add_14_36_groupi_g52789 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_223), .y(csa_tree_add_14_36_groupi_n_340));
nor2 csa_tree_add_14_36_groupi_g52790 (.a(csa_tree_add_14_36_groupi_n_255), .b(csa_tree_add_14_36_groupi_n_204), .y(csa_tree_add_14_36_groupi_n_339));
nand2 csa_tree_add_14_36_groupi_g52791 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_287), .y(csa_tree_add_14_36_groupi_n_338));
nand2 csa_tree_add_14_36_groupi_g52792 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_304), .y(csa_tree_add_14_36_groupi_n_337));
nand2 csa_tree_add_14_36_groupi_g52793 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_288), .y(csa_tree_add_14_36_groupi_n_336));
nand2 csa_tree_add_14_36_groupi_g52794 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_307), .y(csa_tree_add_14_36_groupi_n_335));
nand2 csa_tree_add_14_36_groupi_g52795 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_289), .y(csa_tree_add_14_36_groupi_n_334));
nand2 csa_tree_add_14_36_groupi_g52796 (.a(csa_tree_add_14_36_groupi_n_148), .b(a_0), .y(csa_tree_add_14_36_groupi_n_333));
nand2 csa_tree_add_14_36_groupi_g52797 (.a(csa_tree_add_14_36_groupi_n_146), .b(a_0), .y(csa_tree_add_14_36_groupi_n_332));
nand2 csa_tree_add_14_36_groupi_g52798 (.a(csa_tree_add_14_36_groupi_n_150), .b(a_0), .y(csa_tree_add_14_36_groupi_n_331));
nand2 csa_tree_add_14_36_groupi_g52799 (.a(csa_tree_add_14_36_groupi_n_144), .b(a_0), .y(csa_tree_add_14_36_groupi_n_330));
nand2 csa_tree_add_14_36_groupi_g52800 (.a(csa_tree_add_14_36_groupi_n_257), .b(a_0), .y(csa_tree_add_14_36_groupi_n_329));
nand2 csa_tree_add_14_36_groupi_g52801 (.a(csa_tree_add_14_36_groupi_n_148), .b(b_7), .y(csa_tree_add_14_36_groupi_n_328));
nand2 csa_tree_add_14_36_groupi_g52802 (.a(csa_tree_add_14_36_groupi_n_144), .b(b_13), .y(csa_tree_add_14_36_groupi_n_327));
nand2 csa_tree_add_14_36_groupi_g52803 (.a(csa_tree_add_14_36_groupi_n_257), .b(b_11), .y(csa_tree_add_14_36_groupi_n_326));
nand2 csa_tree_add_14_36_groupi_g52804 (.a(csa_tree_add_14_36_groupi_n_150), .b(b_3), .y(csa_tree_add_14_36_groupi_n_325));
nand2 csa_tree_add_14_36_groupi_g52805 (.a(csa_tree_add_14_36_groupi_n_146), .b(b_5), .y(csa_tree_add_14_36_groupi_n_324));
nand2 csa_tree_add_14_36_groupi_g52806 (.a(csa_tree_add_14_36_groupi_n_254), .b(a_0), .y(csa_tree_add_14_36_groupi_n_323));
nand2 csa_tree_add_14_36_groupi_g52807 (.a(n_2583), .b(a_0), .y(csa_tree_add_14_36_groupi_n_322));
nor2 csa_tree_add_14_36_groupi_g52808 (.a(csa_tree_add_14_36_groupi_n_259), .b(csa_tree_add_14_36_groupi_n_110), .y(csa_tree_add_14_36_groupi_n_321));
nor2 csa_tree_add_14_36_groupi_g52809 (.a(csa_tree_add_14_36_groupi_n_255), .b(csa_tree_add_14_36_groupi_n_236), .y(csa_tree_add_14_36_groupi_n_320));
nand2 csa_tree_add_14_36_groupi_g52810 (.a(csa_tree_add_14_36_groupi_n_254), .b(b_9), .y(csa_tree_add_14_36_groupi_n_319));
nand2 csa_tree_add_14_36_groupi_g52811 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_306), .y(csa_tree_add_14_36_groupi_n_318));
nand2 csa_tree_add_14_36_groupi_g52812 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_305), .y(csa_tree_add_14_36_groupi_n_317));
xor2 csa_tree_add_14_36_groupi_g52813 (.a(csa_tree_add_14_36_groupi_n_98), .b(b_1), .y(csa_tree_add_14_36_groupi_n_316));
nand2 csa_tree_add_14_36_groupi_g52814 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_290), .y(csa_tree_add_14_36_groupi_n_409));
nand2 csa_tree_add_14_36_groupi_g52815 (.a(n_2583), .b(b_15), .y(csa_tree_add_14_36_groupi_n_408));
nor2 csa_tree_add_14_36_groupi_g52816 (.a(csa_tree_add_14_36_groupi_n_254), .b(csa_tree_add_14_36_groupi_n_293), .y(csa_tree_add_14_36_groupi_n_407));
nor2 csa_tree_add_14_36_groupi_g52817 (.a(n_2583), .b(csa_tree_add_14_36_groupi_n_291), .y(csa_tree_add_14_36_groupi_n_404));
inv csa_tree_add_14_36_groupi_g52823 (.a(csa_tree_add_14_36_groupi_n_238), .y(csa_tree_add_14_36_groupi_n_315));
inv csa_tree_add_14_36_groupi_g52824 (.a(csa_tree_add_14_36_groupi_n_2033), .y(csa_tree_add_14_36_groupi_n_298));
inv csa_tree_add_14_36_groupi_g52825 (.a(csa_tree_add_14_36_groupi_n_2027), .y(csa_tree_add_14_36_groupi_n_295));
inv csa_tree_add_14_36_groupi_g52826 (.a(csa_tree_add_14_36_groupi_n_268), .y(csa_tree_add_14_36_groupi_n_269));
inv csa_tree_add_14_36_groupi_g52827 (.a(csa_tree_add_14_36_groupi_n_2028), .y(csa_tree_add_14_36_groupi_n_264));
inv csa_tree_add_14_36_groupi_g52828 (.a(csa_tree_add_14_36_groupi_n_2158), .y(csa_tree_add_14_36_groupi_n_263));
inv csa_tree_add_14_36_groupi_g52829 (.a(csa_tree_add_14_36_groupi_n_2155), .y(csa_tree_add_14_36_groupi_n_262));
inv csa_tree_add_14_36_groupi_g52830 (.a(csa_tree_add_14_36_groupi_n_2034), .y(csa_tree_add_14_36_groupi_n_261));
inv csa_tree_add_14_36_groupi_g52831 (.a(csa_tree_add_14_36_groupi_n_2035), .y(csa_tree_add_14_36_groupi_n_260));
inv csa_tree_add_14_36_groupi_g52834 (.a(csa_tree_add_14_36_groupi_n_255), .y(csa_tree_add_14_36_groupi_n_254));
nor2 csa_tree_add_14_36_groupi_g52835 (.a(csa_tree_add_14_36_groupi_n_124), .b(csa_tree_add_14_36_groupi_n_60), .y(csa_tree_add_14_36_groupi_n_253));
xor2 csa_tree_add_14_36_groupi_g52836 (.a(a_0), .b(b_5), .y(csa_tree_add_14_36_groupi_n_252));
nor2 csa_tree_add_14_36_groupi_g52837 (.a(csa_tree_add_14_36_groupi_n_127), .b(csa_tree_add_14_36_groupi_n_88), .y(csa_tree_add_14_36_groupi_n_251));
nand2 csa_tree_add_14_36_groupi_g52838 (.a(n_2616), .b(csa_tree_add_14_36_groupi_n_92), .y(csa_tree_add_14_36_groupi_n_250));
nor2 csa_tree_add_14_36_groupi_g52839 (.a(n_2616), .b(csa_tree_add_14_36_groupi_n_110), .y(csa_tree_add_14_36_groupi_n_249));
nand2 csa_tree_add_14_36_groupi_g52840 (.a(csa_tree_add_14_36_groupi_n_127), .b(csa_tree_add_14_36_groupi_n_91), .y(csa_tree_add_14_36_groupi_n_248));
nand2 csa_tree_add_14_36_groupi_g52841 (.a(csa_tree_add_14_36_groupi_n_125), .b(b_13), .y(csa_tree_add_14_36_groupi_n_247));
nand2 csa_tree_add_14_36_groupi_g52842 (.a(csa_tree_add_14_36_groupi_n_122), .b(b_5), .y(csa_tree_add_14_36_groupi_n_246));
nand2 csa_tree_add_14_36_groupi_g52843 (.a(csa_tree_add_14_36_groupi_n_120), .b(b_11), .y(csa_tree_add_14_36_groupi_n_245));
nor2 csa_tree_add_14_36_groupi_g52845 (.a(csa_tree_add_14_36_groupi_n_119), .b(csa_tree_add_14_36_groupi_n_59), .y(csa_tree_add_14_36_groupi_n_243));
nor2 csa_tree_add_14_36_groupi_g52846 (.a(csa_tree_add_14_36_groupi_n_123), .b(csa_tree_add_14_36_groupi_n_74), .y(csa_tree_add_14_36_groupi_n_242));
nor2 csa_tree_add_14_36_groupi_g52847 (.a(csa_tree_add_14_36_groupi_n_118), .b(b_1), .y(csa_tree_add_14_36_groupi_n_241));
nor2 csa_tree_add_14_36_groupi_g52849 (.a(csa_tree_add_14_36_groupi_n_113), .b(n_2445), .y(csa_tree_add_14_36_groupi_n_240));
nand2 csa_tree_add_14_36_groupi_g52850 (.a(csa_tree_add_14_36_groupi_n_98), .b(b_1), .y(csa_tree_add_14_36_groupi_n_239));
nor2 csa_tree_add_14_36_groupi_g52851 (.a(csa_tree_add_14_36_groupi_n_98), .b(b_1), .y(csa_tree_add_14_36_groupi_n_238));
nand2 csa_tree_add_14_36_groupi_g52852 (.a(csa_tree_add_14_36_groupi_n_97), .b(csa_tree_add_14_36_groupi_n_76), .y(csa_tree_add_14_36_groupi_n_237));
xor2 csa_tree_add_14_36_groupi_g52853 (.a(csa_tree_add_14_36_groupi_n_74), .b(a_3), .y(csa_tree_add_14_36_groupi_n_236));
xor2 csa_tree_add_14_36_groupi_g52854 (.a(csa_tree_add_14_36_groupi_n_57), .b(a_0), .y(csa_tree_add_14_36_groupi_n_235));
xor2 csa_tree_add_14_36_groupi_g52855 (.a(a_0), .b(b_9), .y(csa_tree_add_14_36_groupi_n_234));
xor2 csa_tree_add_14_36_groupi_g52858 (.a(b_5), .b(b_4), .y(csa_tree_add_14_36_groupi_n_231));
xor2 csa_tree_add_14_36_groupi_g52859 (.a(b_3), .b(b_2), .y(csa_tree_add_14_36_groupi_n_230));
nor2 csa_tree_add_14_36_groupi_g52862 (.a(csa_tree_add_14_36_groupi_n_2250), .b(csa_tree_add_14_36_groupi_n_2240), .y(csa_tree_add_14_36_groupi_n_313));
xor2 csa_tree_add_14_36_groupi_g52863 (.a(a_1), .b(b_11), .y(csa_tree_add_14_36_groupi_n_312));
xor2 csa_tree_add_14_36_groupi_g52864 (.a(a_4), .b(b_11), .y(csa_tree_add_14_36_groupi_n_311));
nor2 csa_tree_add_14_36_groupi_g52865 (.a(csa_tree_add_14_36_groupi_n_100), .b(csa_tree_add_14_36_groupi_n_134), .y(csa_tree_add_14_36_groupi_n_310));
xor2 csa_tree_add_14_36_groupi_g52866 (.a(a_14), .b(b_5), .y(csa_tree_add_14_36_groupi_n_309));
xor2 csa_tree_add_14_36_groupi_g52867 (.a(a_7), .b(b_15), .y(csa_tree_add_14_36_groupi_n_308));
xor2 csa_tree_add_14_36_groupi_g52868 (.a(a_4), .b(b_15), .y(csa_tree_add_14_36_groupi_n_307));
xor2 csa_tree_add_14_36_groupi_g52869 (.a(a_15), .b(b_15), .y(csa_tree_add_14_36_groupi_n_306));
xor2 csa_tree_add_14_36_groupi_g52870 (.a(a_12), .b(b_15), .y(csa_tree_add_14_36_groupi_n_305));
xor2 csa_tree_add_14_36_groupi_g52871 (.a(a_14), .b(b_15), .y(csa_tree_add_14_36_groupi_n_304));
xor2 csa_tree_add_14_36_groupi_g52872 (.a(a_3), .b(b_15), .y(csa_tree_add_14_36_groupi_n_303));
xor2 csa_tree_add_14_36_groupi_g52873 (.a(a_2), .b(b_15), .y(csa_tree_add_14_36_groupi_n_302));
xor2 csa_tree_add_14_36_groupi_g52874 (.a(a_13), .b(b_15), .y(csa_tree_add_14_36_groupi_n_301));
xor2 csa_tree_add_14_36_groupi_g52875 (.a(a_6), .b(b_15), .y(csa_tree_add_14_36_groupi_n_300));
xor2 csa_tree_add_14_36_groupi_g52876 (.a(a_10), .b(b_5), .y(csa_tree_add_14_36_groupi_n_299));
xor2 csa_tree_add_14_36_groupi_g52878 (.a(a_5), .b(b_9), .y(csa_tree_add_14_36_groupi_n_297));
xor2 csa_tree_add_14_36_groupi_g52879 (.a(a_10), .b(b_3), .y(csa_tree_add_14_36_groupi_n_296));
xor2 csa_tree_add_14_36_groupi_g52882 (.a(a_6), .b(b_5), .y(csa_tree_add_14_36_groupi_n_294));
xor2 csa_tree_add_14_36_groupi_g52883 (.a(csa_tree_add_14_36_groupi_n_74), .b(b_8), .y(csa_tree_add_14_36_groupi_n_293));
nand2 csa_tree_add_14_36_groupi_g52884 (.a(n_2537), .b(b_15), .y(csa_tree_add_14_36_groupi_n_292));
xor2 csa_tree_add_14_36_groupi_g52885 (.a(csa_tree_add_14_36_groupi_n_57), .b(b_14), .y(csa_tree_add_14_36_groupi_n_291));
xor2 csa_tree_add_14_36_groupi_g52886 (.a(n_133), .b(n_147), .y(csa_tree_add_14_36_groupi_n_228));
xor2 csa_tree_add_14_36_groupi_g52887 (.a(n_151), .b(n_125), .y(csa_tree_add_14_36_groupi_n_227));
xor2 csa_tree_add_14_36_groupi_g52888 (.a(a_11), .b(b_15), .y(csa_tree_add_14_36_groupi_n_290));
xor2 csa_tree_add_14_36_groupi_g52889 (.a(a_8), .b(b_15), .y(csa_tree_add_14_36_groupi_n_289));
xor2 csa_tree_add_14_36_groupi_g52890 (.a(a_5), .b(b_15), .y(csa_tree_add_14_36_groupi_n_288));
xor2 csa_tree_add_14_36_groupi_g52891 (.a(a_9), .b(b_15), .y(csa_tree_add_14_36_groupi_n_287));
xor2 csa_tree_add_14_36_groupi_g52892 (.a(a_8), .b(b_9), .y(csa_tree_add_14_36_groupi_n_286));
xor2 csa_tree_add_14_36_groupi_g52893 (.a(a_11), .b(b_3), .y(csa_tree_add_14_36_groupi_n_285));
xor2 csa_tree_add_14_36_groupi_g52894 (.a(a_15), .b(b_9), .y(csa_tree_add_14_36_groupi_n_284));
xor2 csa_tree_add_14_36_groupi_g52895 (.a(a_6), .b(b_1), .y(csa_tree_add_14_36_groupi_n_283));
xor2 csa_tree_add_14_36_groupi_g52896 (.a(a_5), .b(b_5), .y(csa_tree_add_14_36_groupi_n_282));
xor2 csa_tree_add_14_36_groupi_g52897 (.a(a_14), .b(b_11), .y(csa_tree_add_14_36_groupi_n_281));
xor2 csa_tree_add_14_36_groupi_g52898 (.a(a_10), .b(b_11), .y(csa_tree_add_14_36_groupi_n_280));
xor2 csa_tree_add_14_36_groupi_g52899 (.a(a_2), .b(b_3), .y(csa_tree_add_14_36_groupi_n_279));
xor2 csa_tree_add_14_36_groupi_g52900 (.a(a_14), .b(b_1), .y(csa_tree_add_14_36_groupi_n_278));
xor2 csa_tree_add_14_36_groupi_g52901 (.a(a_3), .b(b_5), .y(csa_tree_add_14_36_groupi_n_277));
xor2 csa_tree_add_14_36_groupi_g52902 (.a(a_8), .b(b_3), .y(csa_tree_add_14_36_groupi_n_276));
xor2 csa_tree_add_14_36_groupi_g52903 (.a(a_13), .b(b_11), .y(csa_tree_add_14_36_groupi_n_275));
xor2 csa_tree_add_14_36_groupi_g52904 (.a(a_12), .b(b_1), .y(csa_tree_add_14_36_groupi_n_274));
xor2 csa_tree_add_14_36_groupi_g52905 (.a(a_9), .b(b_3), .y(csa_tree_add_14_36_groupi_n_273));
xor2 csa_tree_add_14_36_groupi_g52906 (.a(a_5), .b(b_3), .y(csa_tree_add_14_36_groupi_n_272));
xor2 csa_tree_add_14_36_groupi_g52907 (.a(a_6), .b(b_9), .y(csa_tree_add_14_36_groupi_n_271));
xor2 csa_tree_add_14_36_groupi_g52908 (.a(a_13), .b(b_1), .y(csa_tree_add_14_36_groupi_n_270));
xor2 csa_tree_add_14_36_groupi_g52909 (.a(a_10), .b(b_9), .y(csa_tree_add_14_36_groupi_n_268));
xor2 csa_tree_add_14_36_groupi_g52910 (.a(a_4), .b(b_5), .y(csa_tree_add_14_36_groupi_n_267));
xor2 csa_tree_add_14_36_groupi_g52911 (.a(a_8), .b(b_5), .y(csa_tree_add_14_36_groupi_n_266));
xor2 csa_tree_add_14_36_groupi_g52912 (.a(a_1), .b(b_9), .y(csa_tree_add_14_36_groupi_n_265));
xor2 csa_tree_add_14_36_groupi_g52920 (.a(b_10), .b(b_9), .y(csa_tree_add_14_36_groupi_n_257));
nand2 csa_tree_add_14_36_groupi_g52921 (.a(csa_tree_add_14_36_groupi_n_127), .b(csa_tree_add_14_36_groupi_n_128), .y(csa_tree_add_14_36_groupi_n_255));
inv csa_tree_add_14_36_groupi_g52923 (.a(csa_tree_add_14_36_groupi_n_148), .y(csa_tree_add_14_36_groupi_n_147));
xor2 csa_tree_add_14_36_groupi_g52926 (.a(a_0), .b(b_7), .y(csa_tree_add_14_36_groupi_n_142));
xor2 csa_tree_add_14_36_groupi_g52927 (.a(a_0), .b(b_3), .y(csa_tree_add_14_36_groupi_n_141));
xor2 csa_tree_add_14_36_groupi_g52928 (.a(a_0), .b(b_11), .y(csa_tree_add_14_36_groupi_n_140));
xor2 csa_tree_add_14_36_groupi_g52929 (.a(a_0), .b(b_13), .y(csa_tree_add_14_36_groupi_n_139));
xor2 csa_tree_add_14_36_groupi_g52930 (.a(a_12), .b(b_3), .y(csa_tree_add_14_36_groupi_n_226));
xor2 csa_tree_add_14_36_groupi_g52931 (.a(a_4), .b(b_3), .y(csa_tree_add_14_36_groupi_n_225));
xor2 csa_tree_add_14_36_groupi_g52932 (.a(a_12), .b(b_5), .y(csa_tree_add_14_36_groupi_n_224));
xor2 csa_tree_add_14_36_groupi_g52933 (.a(a_12), .b(b_9), .y(csa_tree_add_14_36_groupi_n_223));
xor2 csa_tree_add_14_36_groupi_g52934 (.a(a_4), .b(b_1), .y(csa_tree_add_14_36_groupi_n_222));
xor2 csa_tree_add_14_36_groupi_g52935 (.a(a_13), .b(b_5), .y(csa_tree_add_14_36_groupi_n_221));
xor2 csa_tree_add_14_36_groupi_g52936 (.a(a_7), .b(b_9), .y(csa_tree_add_14_36_groupi_n_220));
xor2 csa_tree_add_14_36_groupi_g52937 (.a(a_11), .b(b_1), .y(csa_tree_add_14_36_groupi_n_219));
xor2 csa_tree_add_14_36_groupi_g52938 (.a(a_14), .b(b_3), .y(csa_tree_add_14_36_groupi_n_218));
xor2 csa_tree_add_14_36_groupi_g52939 (.a(a_3), .b(b_3), .y(csa_tree_add_14_36_groupi_n_217));
xor2 csa_tree_add_14_36_groupi_g52940 (.a(a_4), .b(b_9), .y(csa_tree_add_14_36_groupi_n_216));
xor2 csa_tree_add_14_36_groupi_g52941 (.a(a_2), .b(b_1), .y(csa_tree_add_14_36_groupi_n_215));
xor2 csa_tree_add_14_36_groupi_g52942 (.a(a_12), .b(b_11), .y(csa_tree_add_14_36_groupi_n_214));
xor2 csa_tree_add_14_36_groupi_g52943 (.a(a_11), .b(b_9), .y(csa_tree_add_14_36_groupi_n_213));
xor2 csa_tree_add_14_36_groupi_g52944 (.a(a_9), .b(b_11), .y(csa_tree_add_14_36_groupi_n_212));
xor2 csa_tree_add_14_36_groupi_g52945 (.a(n_129), .b(n_127), .y(csa_tree_add_14_36_groupi_n_138));
xor2 csa_tree_add_14_36_groupi_g52946 (.a(a_15), .b(b_1), .y(csa_tree_add_14_36_groupi_n_211));
xor2 csa_tree_add_14_36_groupi_g52947 (.a(a_5), .b(b_1), .y(csa_tree_add_14_36_groupi_n_210));
xor2 csa_tree_add_14_36_groupi_g52948 (.a(a_11), .b(b_11), .y(csa_tree_add_14_36_groupi_n_209));
xor2 csa_tree_add_14_36_groupi_g52949 (.a(a_8), .b(b_11), .y(csa_tree_add_14_36_groupi_n_208));
xor2 csa_tree_add_14_36_groupi_g52950 (.a(a_7), .b(b_3), .y(csa_tree_add_14_36_groupi_n_207));
xor2 csa_tree_add_14_36_groupi_g52951 (.a(a_6), .b(b_3), .y(csa_tree_add_14_36_groupi_n_206));
xor2 csa_tree_add_14_36_groupi_g52952 (.a(a_1), .b(b_3), .y(csa_tree_add_14_36_groupi_n_205));
xor2 csa_tree_add_14_36_groupi_g52953 (.a(csa_tree_add_14_36_groupi_n_74), .b(a_9), .y(csa_tree_add_14_36_groupi_n_204));
xor2 csa_tree_add_14_36_groupi_g52954 (.a(a_1), .b(b_1), .y(csa_tree_add_14_36_groupi_n_203));
xor2 csa_tree_add_14_36_groupi_g52955 (.a(a_2), .b(b_11), .y(csa_tree_add_14_36_groupi_n_202));
xor2 csa_tree_add_14_36_groupi_g52956 (.a(a_2), .b(b_5), .y(csa_tree_add_14_36_groupi_n_201));
xor2 csa_tree_add_14_36_groupi_g52957 (.a(a_9), .b(b_5), .y(csa_tree_add_14_36_groupi_n_200));
xor2 csa_tree_add_14_36_groupi_g52958 (.a(n_131), .b(n_149), .y(csa_tree_add_14_36_groupi_n_137));
xor2 csa_tree_add_14_36_groupi_g52959 (.a(a_11), .b(b_5), .y(csa_tree_add_14_36_groupi_n_199));
xor2 csa_tree_add_14_36_groupi_g52960 (.a(a_13), .b(b_3), .y(csa_tree_add_14_36_groupi_n_198));
xor2 csa_tree_add_14_36_groupi_g52961 (.a(n_137), .b(n_145), .y(csa_tree_add_14_36_groupi_n_136));
xor2 csa_tree_add_14_36_groupi_g52962 (.a(a_6), .b(b_11), .y(csa_tree_add_14_36_groupi_n_197));
xor2 csa_tree_add_14_36_groupi_g52963 (.a(a_3), .b(b_11), .y(csa_tree_add_14_36_groupi_n_196));
xor2 csa_tree_add_14_36_groupi_g52964 (.a(a_7), .b(b_5), .y(csa_tree_add_14_36_groupi_n_195));
xor2 csa_tree_add_14_36_groupi_g52965 (.a(a_5), .b(b_11), .y(csa_tree_add_14_36_groupi_n_194));
xor2 csa_tree_add_14_36_groupi_g52966 (.a(a_7), .b(b_11), .y(csa_tree_add_14_36_groupi_n_193));
xor2 csa_tree_add_14_36_groupi_g52967 (.a(a_15), .b(b_5), .y(csa_tree_add_14_36_groupi_n_192));
xor2 csa_tree_add_14_36_groupi_g52968 (.a(a_13), .b(b_9), .y(csa_tree_add_14_36_groupi_n_191));
xor2 csa_tree_add_14_36_groupi_g52969 (.a(n_141), .b(n_139), .y(csa_tree_add_14_36_groupi_n_135));
xor2 csa_tree_add_14_36_groupi_g52970 (.a(a_15), .b(b_3), .y(csa_tree_add_14_36_groupi_n_190));
xor2 csa_tree_add_14_36_groupi_g52971 (.a(a_15), .b(b_11), .y(csa_tree_add_14_36_groupi_n_189));
xor2 csa_tree_add_14_36_groupi_g52972 (.a(a_9), .b(b_1), .y(csa_tree_add_14_36_groupi_n_188));
xor2 csa_tree_add_14_36_groupi_g52973 (.a(a_1), .b(b_5), .y(csa_tree_add_14_36_groupi_n_187));
xor2 csa_tree_add_14_36_groupi_g52974 (.a(a_3), .b(b_1), .y(csa_tree_add_14_36_groupi_n_186));
xor2 csa_tree_add_14_36_groupi_g52975 (.a(a_10), .b(b_1), .y(csa_tree_add_14_36_groupi_n_185));
xor2 csa_tree_add_14_36_groupi_g52976 (.a(a_14), .b(b_9), .y(csa_tree_add_14_36_groupi_n_184));
xor2 csa_tree_add_14_36_groupi_g52977 (.a(a_7), .b(b_1), .y(csa_tree_add_14_36_groupi_n_183));
xor2 csa_tree_add_14_36_groupi_g52978 (.a(a_5), .b(b_13), .y(csa_tree_add_14_36_groupi_n_182));
xor2 csa_tree_add_14_36_groupi_g52979 (.a(a_6), .b(b_7), .y(csa_tree_add_14_36_groupi_n_181));
xor2 csa_tree_add_14_36_groupi_g52980 (.a(a_2), .b(b_7), .y(csa_tree_add_14_36_groupi_n_180));
xor2 csa_tree_add_14_36_groupi_g52981 (.a(a_6), .b(b_13), .y(csa_tree_add_14_36_groupi_n_179));
xor2 csa_tree_add_14_36_groupi_g52982 (.a(a_5), .b(b_7), .y(csa_tree_add_14_36_groupi_n_178));
xor2 csa_tree_add_14_36_groupi_g52983 (.a(a_3), .b(b_13), .y(csa_tree_add_14_36_groupi_n_177));
xor2 csa_tree_add_14_36_groupi_g52984 (.a(a_4), .b(b_13), .y(csa_tree_add_14_36_groupi_n_176));
xor2 csa_tree_add_14_36_groupi_g52985 (.a(a_1), .b(b_13), .y(csa_tree_add_14_36_groupi_n_175));
xor2 csa_tree_add_14_36_groupi_g52986 (.a(a_12), .b(b_7), .y(csa_tree_add_14_36_groupi_n_174));
xor2 csa_tree_add_14_36_groupi_g52987 (.a(a_11), .b(b_7), .y(csa_tree_add_14_36_groupi_n_173));
xor2 csa_tree_add_14_36_groupi_g52988 (.a(a_8), .b(b_7), .y(csa_tree_add_14_36_groupi_n_172));
xor2 csa_tree_add_14_36_groupi_g52989 (.a(a_7), .b(b_13), .y(csa_tree_add_14_36_groupi_n_171));
xor2 csa_tree_add_14_36_groupi_g52990 (.a(a_8), .b(b_1), .y(csa_tree_add_14_36_groupi_n_170));
xor2 csa_tree_add_14_36_groupi_g52991 (.a(a_13), .b(b_13), .y(csa_tree_add_14_36_groupi_n_169));
xor2 csa_tree_add_14_36_groupi_g52992 (.a(a_8), .b(b_13), .y(csa_tree_add_14_36_groupi_n_168));
xor2 csa_tree_add_14_36_groupi_g52993 (.a(a_15), .b(b_13), .y(csa_tree_add_14_36_groupi_n_167));
xor2 csa_tree_add_14_36_groupi_g52994 (.a(a_11), .b(b_13), .y(csa_tree_add_14_36_groupi_n_166));
xor2 csa_tree_add_14_36_groupi_g52995 (.a(a_14), .b(b_13), .y(csa_tree_add_14_36_groupi_n_165));
xor2 csa_tree_add_14_36_groupi_g52996 (.a(a_4), .b(b_7), .y(csa_tree_add_14_36_groupi_n_164));
xor2 csa_tree_add_14_36_groupi_g52997 (.a(csa_tree_add_14_36_groupi_n_74), .b(a_2), .y(csa_tree_add_14_36_groupi_n_163));
xor2 csa_tree_add_14_36_groupi_g52998 (.a(a_3), .b(b_7), .y(csa_tree_add_14_36_groupi_n_162));
xor2 csa_tree_add_14_36_groupi_g52999 (.a(a_14), .b(b_7), .y(csa_tree_add_14_36_groupi_n_161));
xor2 csa_tree_add_14_36_groupi_g53000 (.a(a_15), .b(b_7), .y(csa_tree_add_14_36_groupi_n_160));
xor2 csa_tree_add_14_36_groupi_g53001 (.a(a_10), .b(b_13), .y(csa_tree_add_14_36_groupi_n_159));
xor2 csa_tree_add_14_36_groupi_g53002 (.a(a_13), .b(b_7), .y(csa_tree_add_14_36_groupi_n_158));
xor2 csa_tree_add_14_36_groupi_g53003 (.a(a_7), .b(b_7), .y(csa_tree_add_14_36_groupi_n_157));
xor2 csa_tree_add_14_36_groupi_g53004 (.a(a_10), .b(b_7), .y(csa_tree_add_14_36_groupi_n_156));
xor2 csa_tree_add_14_36_groupi_g53005 (.a(a_2), .b(b_13), .y(csa_tree_add_14_36_groupi_n_155));
xor2 csa_tree_add_14_36_groupi_g53006 (.a(a_9), .b(b_13), .y(csa_tree_add_14_36_groupi_n_154));
xor2 csa_tree_add_14_36_groupi_g53007 (.a(a_1), .b(b_7), .y(csa_tree_add_14_36_groupi_n_153));
xor2 csa_tree_add_14_36_groupi_g53008 (.a(a_12), .b(b_13), .y(csa_tree_add_14_36_groupi_n_152));
xor2 csa_tree_add_14_36_groupi_g53009 (.a(a_9), .b(b_7), .y(csa_tree_add_14_36_groupi_n_151));
xor2 csa_tree_add_14_36_groupi_g53010 (.a(b_2), .b(b_1), .y(csa_tree_add_14_36_groupi_n_150));
xor2 csa_tree_add_14_36_groupi_g53011 (.a(b_6), .b(b_5), .y(csa_tree_add_14_36_groupi_n_148));
xor2 csa_tree_add_14_36_groupi_g53012 (.a(b_4), .b(b_3), .y(csa_tree_add_14_36_groupi_n_146));
xor2 csa_tree_add_14_36_groupi_g53013 (.a(b_12), .b(b_11), .y(csa_tree_add_14_36_groupi_n_144));
inv csa_tree_add_14_36_groupi_g53015 (.a(csa_tree_add_14_36_groupi_n_2250), .y(csa_tree_add_14_36_groupi_n_130));
inv csa_tree_add_14_36_groupi_g53016 (.a(csa_tree_add_14_36_groupi_n_129), .y(csa_tree_add_14_36_groupi_n_128));
nand2 csa_tree_add_14_36_groupi_g53018 (.a(a_0), .b(b_12), .y(csa_tree_add_14_36_groupi_n_125));
nor2 csa_tree_add_14_36_groupi_g53019 (.a(a_0), .b(b_12), .y(csa_tree_add_14_36_groupi_n_124));
nor2 csa_tree_add_14_36_groupi_g53020 (.a(a_0), .b(b_10), .y(csa_tree_add_14_36_groupi_n_123));
nand2 csa_tree_add_14_36_groupi_g53021 (.a(a_0), .b(b_4), .y(csa_tree_add_14_36_groupi_n_122));
nor2 csa_tree_add_14_36_groupi_g53022 (.a(a_0), .b(b_6), .y(csa_tree_add_14_36_groupi_n_121));
nand2 csa_tree_add_14_36_groupi_g53023 (.a(a_0), .b(b_10), .y(csa_tree_add_14_36_groupi_n_120));
nor2 csa_tree_add_14_36_groupi_g53024 (.a(a_0), .b(b_4), .y(csa_tree_add_14_36_groupi_n_119));
nor2 csa_tree_add_14_36_groupi_g53025 (.a(csa_tree_add_14_36_groupi_n_76), .b(csa_tree_add_14_36_groupi_n_78), .y(csa_tree_add_14_36_groupi_n_118));
nor2 csa_tree_add_14_36_groupi_g53026 (.a(a_0), .b(b_2), .y(csa_tree_add_14_36_groupi_n_117));
nand2 csa_tree_add_14_36_groupi_g53027 (.a(a_4), .b(b_15), .y(csa_tree_add_14_36_groupi_n_116));
nor2 csa_tree_add_14_36_groupi_g53028 (.a(a_10), .b(b_15), .y(csa_tree_add_14_36_groupi_n_134));
nand2 csa_tree_add_14_36_groupi_g53030 (.a(a_15), .b(b_15), .y(csa_tree_add_14_36_groupi_n_115));
nand2 csa_tree_add_14_36_groupi_g53031 (.a(a_6), .b(b_15), .y(csa_tree_add_14_36_groupi_n_114));
nor2 csa_tree_add_14_36_groupi_g53035 (.a(b_8), .b(b_7), .y(csa_tree_add_14_36_groupi_n_129));
nand2 csa_tree_add_14_36_groupi_g53036 (.a(b_8), .b(b_7), .y(csa_tree_add_14_36_groupi_n_127));
inv csa_tree_add_14_36_groupi_g53037 (.a(n_2508), .y(csa_tree_add_14_36_groupi_n_112));
inv csa_tree_add_14_36_groupi_g53038 (.a(n_2516), .y(csa_tree_add_14_36_groupi_n_109));
inv csa_tree_add_14_36_groupi_g53039 (.a(n_2521), .y(csa_tree_add_14_36_groupi_n_107));
inv csa_tree_add_14_36_groupi_g53040 (.a(csa_tree_add_14_36_groupi_n_103), .y(csa_tree_add_14_36_groupi_n_104));
inv csa_tree_add_14_36_groupi_g53041 (.a(csa_tree_add_14_36_groupi_n_101), .y(csa_tree_add_14_36_groupi_n_102));
inv csa_tree_add_14_36_groupi_g53042 (.a(csa_tree_add_14_36_groupi_n_99), .y(csa_tree_add_14_36_groupi_n_100));
nand2 csa_tree_add_14_36_groupi_g53044 (.a(b_1), .b(b_0), .y(csa_tree_add_14_36_groupi_n_95));
nand2 csa_tree_add_14_36_groupi_g53045 (.a(a_12), .b(b_15), .y(csa_tree_add_14_36_groupi_n_94));
nand2 csa_tree_add_14_36_groupi_g53046 (.a(a_7), .b(b_15), .y(csa_tree_add_14_36_groupi_n_93));
nor2 csa_tree_add_14_36_groupi_g53047 (.a(csa_tree_add_14_36_groupi_n_57), .b(a_0), .y(csa_tree_add_14_36_groupi_n_92));
nor2 csa_tree_add_14_36_groupi_g53048 (.a(csa_tree_add_14_36_groupi_n_74), .b(a_0), .y(csa_tree_add_14_36_groupi_n_91));
nor2 csa_tree_add_14_36_groupi_g53049 (.a(csa_tree_add_14_36_groupi_n_76), .b(csa_tree_add_14_36_groupi_n_77), .y(csa_tree_add_14_36_groupi_n_113));
nand2 csa_tree_add_14_36_groupi_g53051 (.a(a_1), .b(csa_tree_add_14_36_groupi_n_57), .y(csa_tree_add_14_36_groupi_n_110));
nand2 csa_tree_add_14_36_groupi_g53053 (.a(a_13), .b(b_15), .y(csa_tree_add_14_36_groupi_n_90));
nand2 csa_tree_add_14_36_groupi_g53055 (.a(a_14), .b(b_15), .y(csa_tree_add_14_36_groupi_n_89));
nand2 csa_tree_add_14_36_groupi_g53056 (.a(a_3), .b(csa_tree_add_14_36_groupi_n_74), .y(csa_tree_add_14_36_groupi_n_88));
nand2 csa_tree_add_14_36_groupi_g53058 (.a(a_2), .b(b_15), .y(csa_tree_add_14_36_groupi_n_103));
nand2 csa_tree_add_14_36_groupi_g53059 (.a(a_3), .b(b_15), .y(csa_tree_add_14_36_groupi_n_101));
nand2 csa_tree_add_14_36_groupi_g53060 (.a(a_10), .b(b_15), .y(csa_tree_add_14_36_groupi_n_99));
nand2 csa_tree_add_14_36_groupi_g53061 (.a(a_1), .b(b_15), .y(csa_tree_add_14_36_groupi_n_98));
nor2 csa_tree_add_14_36_groupi_g53062 (.a(n_2445), .b(b_0), .y(csa_tree_add_14_36_groupi_n_97));
inv csa_tree_add_14_36_groupi_g53063 (.a(csa_tree_add_14_36_groupi_n_2309), .y(csa_tree_add_14_36_groupi_n_87));
inv csa_tree_add_14_36_groupi_g53064 (.a(n_121), .y(csa_tree_add_14_36_groupi_n_86));
inv csa_tree_add_14_36_groupi_g53065 (.a(csa_tree_add_14_36_groupi_n_2311), .y(csa_tree_add_14_36_groupi_n_85));
inv csa_tree_add_14_36_groupi_g53066 (.a(csa_tree_add_14_36_groupi_n_2315), .y(csa_tree_add_14_36_groupi_n_84));
inv csa_tree_add_14_36_groupi_g53067 (.a(n_75), .y(csa_tree_add_14_36_groupi_n_83));
inv csa_tree_add_14_36_groupi_g53068 (.a(n_82), .y(csa_tree_add_14_36_groupi_n_82));
inv csa_tree_add_14_36_groupi_g53069 (.a(n_153), .y(csa_tree_add_14_36_groupi_n_81));
inv csa_tree_add_14_36_groupi_g53070 (.a(n_125), .y(csa_tree_add_14_36_groupi_n_80));
inv csa_tree_add_14_36_groupi_g53071 (.a(b_6), .y(csa_tree_add_14_36_groupi_n_79));
inv csa_tree_add_14_36_groupi_g53072 (.a(b_2), .y(csa_tree_add_14_36_groupi_n_78));
inv csa_tree_add_14_36_groupi_g53073 (.a(b_0), .y(csa_tree_add_14_36_groupi_n_77));
inv csa_tree_add_14_36_groupi_g53074 (.a(a_0), .y(csa_tree_add_14_36_groupi_n_76));
inv csa_tree_add_14_36_groupi_g53075 (.a(b_7), .y(csa_tree_add_14_36_groupi_n_75));
inv csa_tree_add_14_36_groupi_g53076 (.a(b_9), .y(csa_tree_add_14_36_groupi_n_74));
inv csa_tree_add_14_36_groupi_g53077 (.a(n_78), .y(csa_tree_add_14_36_groupi_n_73));
inv csa_tree_add_14_36_groupi_g53078 (.a(n_123), .y(csa_tree_add_14_36_groupi_n_72));
inv csa_tree_add_14_36_groupi_g53080 (.a(n_159), .y(csa_tree_add_14_36_groupi_n_70));
inv csa_tree_add_14_36_groupi_g53081 (.a(n_80), .y(csa_tree_add_14_36_groupi_n_69));
inv csa_tree_add_14_36_groupi_g53083 (.a(n_76), .y(csa_tree_add_14_36_groupi_n_67));
inv csa_tree_add_14_36_groupi_g53085 (.a(csa_tree_add_14_36_groupi_n_2307), .y(csa_tree_add_14_36_groupi_n_65));
inv csa_tree_add_14_36_groupi_g53086 (.a(csa_tree_add_14_36_groupi_n_2316), .y(csa_tree_add_14_36_groupi_n_64));
inv csa_tree_add_14_36_groupi_g53087 (.a(n_137), .y(csa_tree_add_14_36_groupi_n_63));
inv csa_tree_add_14_36_groupi_g53088 (.a(n_147), .y(csa_tree_add_14_36_groupi_n_62));
inv csa_tree_add_14_36_groupi_g53089 (.a(n_149), .y(csa_tree_add_14_36_groupi_n_61));
inv csa_tree_add_14_36_groupi_g53090 (.a(b_11), .y(csa_tree_add_14_36_groupi_n_60));
inv csa_tree_add_14_36_groupi_g53091 (.a(b_3), .y(csa_tree_add_14_36_groupi_n_59));
inv csa_tree_add_14_36_groupi_g53093 (.a(b_15), .y(csa_tree_add_14_36_groupi_n_57));
inv csa_tree_add_14_36_groupi_g3 (.a(csa_tree_add_14_36_groupi_n_54), .y(csa_tree_add_14_36_groupi_n_53));
nand2 csa_tree_add_14_36_groupi_g2 (.a(csa_tree_add_14_36_groupi_n_1811), .b(n_2488), .y(csa_tree_add_14_36_groupi_n_54));
inv csa_tree_add_14_36_groupi_g53094 (.a(csa_tree_add_14_36_groupi_n_56), .y(csa_tree_add_14_36_groupi_n_52));
nor2 csa_tree_add_14_36_groupi_g53095 (.a(csa_tree_add_14_36_groupi_n_1824), .b(csa_tree_add_14_36_groupi_n_1756), .y(csa_tree_add_14_36_groupi_n_56));
inv csa_tree_add_14_36_groupi_g53096 (.a(csa_tree_add_14_36_groupi_n_51), .y(csa_tree_add_14_36_groupi_n_50));
nand2 csa_tree_add_14_36_groupi_g53097 (.a(csa_tree_add_14_36_groupi_n_1808), .b(csa_tree_add_14_36_groupi_n_1810), .y(csa_tree_add_14_36_groupi_n_51));
inv csa_tree_add_14_36_groupi_g53098 (.a(csa_tree_add_14_36_groupi_n_49), .y(csa_tree_add_14_36_groupi_n_48));
nand2 csa_tree_add_14_36_groupi_g53099 (.a(csa_tree_add_14_36_groupi_n_1569), .b(csa_tree_add_14_36_groupi_n_1728), .y(csa_tree_add_14_36_groupi_n_49));
inv csa_tree_add_14_36_groupi_g53102 (.a(csa_tree_add_14_36_groupi_n_46), .y(csa_tree_add_14_36_groupi_n_45));
nor2 csa_tree_add_14_36_groupi_g53103 (.a(csa_tree_add_14_36_groupi_n_1352), .b(csa_tree_add_14_36_groupi_n_1181), .y(csa_tree_add_14_36_groupi_n_46));
inv csa_tree_add_14_36_groupi_g53104 (.a(csa_tree_add_14_36_groupi_n_44), .y(csa_tree_add_14_36_groupi_n_43));
nand2 csa_tree_add_14_36_groupi_g53105 (.a(csa_tree_add_14_36_groupi_n_1362), .b(csa_tree_add_14_36_groupi_n_1363), .y(csa_tree_add_14_36_groupi_n_44));
inv csa_tree_add_14_36_groupi_g53106 (.a(csa_tree_add_14_36_groupi_n_42), .y(csa_tree_add_14_36_groupi_n_41));
nand2 csa_tree_add_14_36_groupi_g53107 (.a(csa_tree_add_14_36_groupi_n_808), .b(csa_tree_add_14_36_groupi_n_810), .y(csa_tree_add_14_36_groupi_n_42));
dff csa_tree_add_14_36_groupi_retime_s26_6_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_40), .q(csa_tree_add_14_36_groupi_n_2312));
xor2 csa_tree_add_14_36_groupi_g32428 (.a(csa_tree_add_14_36_groupi_n_30), .b(csa_tree_add_14_36_groupi_n_39), .y(csa_tree_add_14_36_groupi_n_40));
xor2 csa_tree_add_14_36_groupi_g32429 (.a(csa_tree_add_14_36_groupi_n_28), .b(csa_tree_add_14_36_groupi_n_36), .y(csa_tree_add_14_36_groupi_n_39));
dff csa_tree_add_14_36_groupi_retime_s20_7_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_37), .q(csa_tree_add_14_36_groupi_n_2308));
dff csa_tree_add_14_36_groupi_retime_s5_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_38), .q(csa_tree_add_14_36_groupi_n_2320));
dff csa_tree_add_14_36_groupi_retime_s26_7_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_33), .q(csa_tree_add_14_36_groupi_n_2311));
dff csa_tree_add_14_36_groupi_retime_s17_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_32), .q(csa_tree_add_14_36_groupi_n_2307));
dff csa_tree_add_14_36_groupi_retime_s2_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_34), .q(csa_tree_add_14_36_groupi_n_2321));
dff csa_tree_add_14_36_groupi_retime_s14_5_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_35), .q(csa_tree_add_14_36_groupi_n_2306));
dff csa_tree_add_14_36_groupi_retime_s23_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_31), .q(csa_tree_add_14_36_groupi_n_2314));
xor2 csa_tree_add_14_36_groupi_g32437 (.a(csa_tree_add_14_36_groupi_n_2281), .b(csa_tree_add_14_36_groupi_n_21), .y(csa_tree_add_14_36_groupi_n_38));
xor2 csa_tree_add_14_36_groupi_g32438 (.a(csa_tree_add_14_36_groupi_n_2286), .b(csa_tree_add_14_36_groupi_n_17), .y(csa_tree_add_14_36_groupi_n_37));
dff csa_tree_add_14_36_groupi_retime_s23_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_29), .q(csa_tree_add_14_36_groupi_n_2309));
xor2 csa_tree_add_14_36_groupi_g32440 (.a(csa_tree_add_14_36_groupi_n_23), .b(csa_tree_add_14_36_groupi_n_24), .y(csa_tree_add_14_36_groupi_n_36));
xor2 csa_tree_add_14_36_groupi_g32441 (.a(csa_tree_add_14_36_groupi_n_20), .b(csa_tree_add_14_36_groupi_n_2278), .y(csa_tree_add_14_36_groupi_n_35));
xor2 csa_tree_add_14_36_groupi_g32442 (.a(csa_tree_add_14_36_groupi_n_2291), .b(n_2623), .y(csa_tree_add_14_36_groupi_n_34));
xor2 csa_tree_add_14_36_groupi_g32443 (.a(csa_tree_add_14_36_groupi_n_2284), .b(csa_tree_add_14_36_groupi_n_19), .y(csa_tree_add_14_36_groupi_n_33));
xor2 csa_tree_add_14_36_groupi_g32444 (.a(csa_tree_add_14_36_groupi_n_2269), .b(csa_tree_add_14_36_groupi_n_18), .y(csa_tree_add_14_36_groupi_n_32));
xor2 csa_tree_add_14_36_groupi_g32445 (.a(csa_tree_add_14_36_groupi_n_2277), .b(csa_tree_add_14_36_groupi_n_25), .y(csa_tree_add_14_36_groupi_n_31));
nand2 csa_tree_add_14_36_groupi_g32446 (.a(csa_tree_add_14_36_groupi_n_26), .b(csa_tree_add_14_36_groupi_n_13), .y(csa_tree_add_14_36_groupi_n_30));
xor2 csa_tree_add_14_36_groupi_g32447 (.a(csa_tree_add_14_36_groupi_n_2292), .b(csa_tree_add_14_36_groupi_n_3), .y(csa_tree_add_14_36_groupi_n_29));
nand2 csa_tree_add_14_36_groupi_g32448 (.a(csa_tree_add_14_36_groupi_n_27), .b(csa_tree_add_14_36_groupi_n_15), .y(csa_tree_add_14_36_groupi_n_28));
dff csa_tree_add_14_36_groupi_retime_s15_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_8), .q(csa_tree_add_14_36_groupi_n_2317));
dff csa_tree_add_14_36_groupi_retime_s26_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_5), .q(csa_tree_add_14_36_groupi_n_2313));
dff csa_tree_add_14_36_groupi_retime_s27_8_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_4), .q(csa_tree_add_14_36_groupi_n_2310));
dff csa_tree_add_14_36_groupi_retime_s8_10_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_9), .q(csa_tree_add_14_36_groupi_n_2303));
dff csa_tree_add_14_36_groupi_retime_s12_2_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_10), .q(csa_tree_add_14_36_groupi_n_2305));
dff csa_tree_add_14_36_groupi_retime_s18_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_7), .q(csa_tree_add_14_36_groupi_n_2316));
nand2 csa_tree_add_14_36_groupi_g32455 (.a(csa_tree_add_14_36_groupi_n_14), .b(csa_tree_add_14_36_groupi_n_2302), .y(csa_tree_add_14_36_groupi_n_27));
nand2 csa_tree_add_14_36_groupi_g32456 (.a(csa_tree_add_14_36_groupi_n_16), .b(csa_tree_add_14_36_groupi_n_2272), .y(csa_tree_add_14_36_groupi_n_26));
xor2 csa_tree_add_14_36_groupi_g32457 (.a(csa_tree_add_14_36_groupi_n_2276), .b(csa_tree_add_14_36_groupi_n_2275), .y(csa_tree_add_14_36_groupi_n_25));
xor2 csa_tree_add_14_36_groupi_g32458 (.a(csa_tree_add_14_36_groupi_n_2297), .b(csa_tree_add_14_36_groupi_n_2298), .y(csa_tree_add_14_36_groupi_n_24));
xor2 csa_tree_add_14_36_groupi_g32459 (.a(n_143), .b(n_135), .y(csa_tree_add_14_36_groupi_n_23));
xor2 csa_tree_add_14_36_groupi_g32461 (.a(csa_tree_add_14_36_groupi_n_2283), .b(csa_tree_add_14_36_groupi_n_2282), .y(csa_tree_add_14_36_groupi_n_21));
xor2 csa_tree_add_14_36_groupi_g32462 (.a(csa_tree_add_14_36_groupi_n_2280), .b(csa_tree_add_14_36_groupi_n_2279), .y(csa_tree_add_14_36_groupi_n_20));
xor2 csa_tree_add_14_36_groupi_g32463 (.a(csa_tree_add_14_36_groupi_n_2285), .b(csa_tree_add_14_36_groupi_n_2300), .y(csa_tree_add_14_36_groupi_n_19));
xor2 csa_tree_add_14_36_groupi_g32464 (.a(csa_tree_add_14_36_groupi_n_2301), .b(csa_tree_add_14_36_groupi_n_2299), .y(csa_tree_add_14_36_groupi_n_18));
xor2 csa_tree_add_14_36_groupi_g32465 (.a(csa_tree_add_14_36_groupi_n_1), .b(csa_tree_add_14_36_groupi_n_2287), .y(csa_tree_add_14_36_groupi_n_17));
inv csa_tree_add_14_36_groupi_g32466 (.a(n_2646), .y(csa_tree_add_14_36_groupi_n_16));
inv csa_tree_add_14_36_groupi_g32467 (.a(csa_tree_add_14_36_groupi_n_11), .y(csa_tree_add_14_36_groupi_n_15));
nand2 csa_tree_add_14_36_groupi_g32468 (.a(n_135), .b(csa_tree_add_14_36_groupi_n_2304), .y(csa_tree_add_14_36_groupi_n_14));
dff csa_tree_add_14_36_groupi_retime_s12_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_2410), .q(csa_tree_add_14_36_groupi_n_2318));
dff csa_tree_add_14_36_groupi_retime_s21_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_2412), .q(csa_tree_add_14_36_groupi_n_2315));
nand2 csa_tree_add_14_36_groupi_g32471 (.a(n_2609), .b(n_2605), .y(csa_tree_add_14_36_groupi_n_13));
nor2 csa_tree_add_14_36_groupi_g32473 (.a(n_135), .b(csa_tree_add_14_36_groupi_n_2304), .y(csa_tree_add_14_36_groupi_n_11));
dff csa_tree_add_14_36_groupi_retime_s8_1_reg (.reset(reset), .ck(clk), .d(csa_tree_add_14_36_groupi_n_2416), .q(csa_tree_add_14_36_groupi_n_2319));
inv csa_tree_add_14_36_groupi_g32475 (.a(csa_tree_add_14_36_groupi_n_6), .y(csa_tree_add_14_36_groupi_n_10));
nand2 csa_tree_add_14_36_groupi_g32476 (.a(csa_tree_add_14_36_groupi_n_2267), .b(csa_tree_add_14_36_groupi_n_2), .y(csa_tree_add_14_36_groupi_n_9));
nand2 csa_tree_add_14_36_groupi_g32477 (.a(csa_tree_add_14_36_groupi_n_2293), .b(csa_tree_add_14_36_groupi_n_2294), .y(csa_tree_add_14_36_groupi_n_8));
nor2 csa_tree_add_14_36_groupi_g32478 (.a(csa_tree_add_14_36_groupi_n_2295), .b(n_2480), .y(csa_tree_add_14_36_groupi_n_7));
nand2 csa_tree_add_14_36_groupi_g32479 (.a(csa_tree_add_14_36_groupi_n_2263), .b(csa_tree_add_14_36_groupi_n_2265), .y(csa_tree_add_14_36_groupi_n_6));
nor2 csa_tree_add_14_36_groupi_g32480 (.a(csa_tree_add_14_36_groupi_n_2270), .b(csa_tree_add_14_36_groupi_n_2271), .y(csa_tree_add_14_36_groupi_n_5));
nand2 csa_tree_add_14_36_groupi_g32481 (.a(csa_tree_add_14_36_groupi_n_2266), .b(csa_tree_add_14_36_groupi_n_0), .y(csa_tree_add_14_36_groupi_n_4));
nand2 csa_tree_add_14_36_groupi_g32482 (.a(csa_tree_add_14_36_groupi_n_2264), .b(csa_tree_add_14_36_groupi_n_2262), .y(csa_tree_add_14_36_groupi_n_3));
inv csa_tree_add_14_36_groupi_g32483 (.a(csa_tree_add_14_36_groupi_n_2268), .y(csa_tree_add_14_36_groupi_n_2));
inv csa_tree_add_14_36_groupi_g32484 (.a(csa_tree_add_14_36_groupi_n_2288), .y(csa_tree_add_14_36_groupi_n_1));
inv csa_tree_add_14_36_groupi_g32485 (.a(csa_tree_add_14_36_groupi_n_2261), .y(csa_tree_add_14_36_groupi_n_0));
nand2 g220 (.a(n_2428), .b(n_2435), .y(n_2436));
inv g226 (.a(n_2427), .y(n_2428));
nor2 g227 (.a(n_2424), .b(n_2426), .y(n_2427));
nor2 g232 (.a(n_2760), .b(csa_tree_add_14_36_groupi_n_1407), .y(n_2424));
inv g233 (.a(n_2425), .y(n_2426));
nand2 g234 (.a(csa_tree_add_14_36_groupi_n_965), .b(csa_tree_add_14_36_groupi_n_1263), .y(n_2425));
nor2 g221 (.a(n_2431), .b(n_2434), .y(n_2435));
nor2 g225 (.a(n_2429), .b(n_2430), .y(n_2431));
nand2 g231 (.a(csa_tree_add_14_36_groupi_n_1204), .b(csa_tree_add_14_36_groupi_n_991), .y(n_2429));
xor2 g229 (.a(csa_tree_add_14_36_groupi_n_1133), .b(csa_tree_add_14_36_groupi_n_1449), .y(n_2430));
nor2 g223 (.a(n_2432), .b(n_2433), .y(n_2434));
xor2 g228 (.a(csa_tree_add_14_36_groupi_n_1087), .b(csa_tree_add_14_36_groupi_n_1048), .y(n_2432));
nand2 g230 (.a(csa_tree_add_14_36_groupi_n_1104), .b(csa_tree_add_14_36_groupi_n_975), .y(n_2433));
nor2 g222 (.a(n_2427), .b(n_2434), .y(n_2437));
inv g224 (.a(n_2431), .y(n_2438));
nand2 g6 (.a(a_0), .b(b_15), .y(n_2440));
inv g2 (.a(b_1), .y(n_2445));
nor2 g15 (.a(n_2450), .b(b_5), .y(n_2451));
nor2 g16 (.a(csa_tree_add_14_36_groupi_n_76), .b(csa_tree_add_14_36_groupi_n_79), .y(n_2450));
nor2 g53108 (.a(n_2659), .b(csa_tree_add_14_36_groupi_n_257), .y(n_2453));
nand2 csa_tree_add_14_36_groupi_g53109 (.a(n_2455), .b(n_2659), .y(n_2457));
inv csa_tree_add_14_36_groupi_g53110 (.a(csa_tree_add_14_36_groupi_n_257), .y(n_2455));
nand2 g9 (.a(n_2458), .b(b_11), .y(n_2459));
inv g10 (.a(n_2453), .y(n_2458));
inv g53112 (.a(n_2460), .y(n_2461));
nor2 g53113 (.a(csa_tree_add_14_36_groupi_n_146), .b(csa_tree_add_14_36_groupi_n_231), .y(n_2460));
nand2 csa_tree_add_14_36_groupi_g53114 (.a(n_2462), .b(csa_tree_add_14_36_groupi_n_231), .y(n_2463));
inv csa_tree_add_14_36_groupi_g53115 (.a(csa_tree_add_14_36_groupi_n_146), .y(n_2462));
nand2 g53116 (.a(n_2464), .b(b_7), .y(n_2465));
nand2 g53117 (.a(b_6), .b(csa_tree_add_14_36_groupi_n_147), .y(n_2464));
nand2 csa_tree_add_14_36_groupi_g53118 (.a(csa_tree_add_14_36_groupi_n_147), .b(n_2466), .y(n_2467));
xor2 csa_tree_add_14_36_groupi_g53119 (.a(b_7), .b(b_6), .y(n_2466));
xor2 g53120 (.a(csa_tree_add_14_36_groupi_n_2306), .b(csa_tree_add_14_36_groupi_n_2256), .y(n_2468));
nand2 csa_tree_add_14_36_groupi_g51282__53121 (.a(n_2469), .b(csa_tree_add_14_36_groupi_n_2256), .y(n_2470));
inv csa_tree_add_14_36_groupi_g53122 (.a(csa_tree_add_14_36_groupi_n_2306), .y(n_2469));
nand2 csa_tree_add_14_36_groupi_g51283__53123 (.a(csa_tree_add_14_36_groupi_n_2306), .b(n_2471), .y(n_2472));
inv csa_tree_add_14_36_groupi_g53124 (.a(csa_tree_add_14_36_groupi_n_2256), .y(n_2471));
nor2 csa_tree_add_14_36_groupi_g51370__53127 (.a(csa_tree_add_14_36_groupi_n_2308), .b(n_2475), .y(n_2476));
inv csa_tree_add_14_36_groupi_g53128 (.a(csa_tree_add_14_36_groupi_n_2208), .y(n_2475));
nor2 csa_tree_add_14_36_groupi_g51361__53129 (.a(n_2477), .b(csa_tree_add_14_36_groupi_n_2208), .y(n_2478));
inv csa_tree_add_14_36_groupi_g53130 (.a(csa_tree_add_14_36_groupi_n_2308), .y(n_2477));
xor2 csa_tree_add_14_36_groupi_g51103__53131 (.a(n_2479), .b(csa_tree_add_14_36_groupi_n_2218), .y(n_2480));
xor2 g53132 (.a(csa_tree_add_14_36_groupi_n_2308), .b(csa_tree_add_14_36_groupi_n_2208), .y(n_2479));
nor2 g22 (.a(n_2482), .b(n_2484), .y(n_2485));
inv g26 (.a(csa_tree_add_14_36_groupi_n_1654), .y(n_2482));
nand2 g24 (.a(csa_tree_add_14_36_groupi_n_1483), .b(n_2483), .y(n_2484));
inv g25 (.a(csa_tree_add_14_36_groupi_n_2249), .y(n_2483));
nand2 g23 (.a(csa_tree_add_14_36_groupi_n_1654), .b(csa_tree_add_14_36_groupi_n_1483), .y(n_2486));
xor2 g53135 (.a(n_2487), .b(csa_tree_add_14_36_groupi_n_2222), .y(n_2488));
xor2 g53136 (.a(csa_tree_add_14_36_groupi_n_2253), .b(csa_tree_add_14_36_groupi_n_2225), .y(n_2487));
nand2 csa_tree_add_14_36_groupi_g51150__53137 (.a(n_2489), .b(csa_tree_add_14_36_groupi_n_2225), .y(n_2490));
inv csa_tree_add_14_36_groupi_g53138 (.a(csa_tree_add_14_36_groupi_n_2253), .y(n_2489));
nand2 csa_tree_add_14_36_groupi_g51152__53139 (.a(csa_tree_add_14_36_groupi_n_2253), .b(n_2491), .y(n_2492));
inv csa_tree_add_14_36_groupi_g53140 (.a(csa_tree_add_14_36_groupi_n_2225), .y(n_2491));
nor2 g53141 (.a(n_2503), .b(n_2504), .y(n_2505));
nand2 g53142 (.a(csa_tree_add_14_36_groupi_n_1871), .b(csa_tree_add_14_36_groupi_n_1834), .y(n_2503));
inv g27 (.a(csa_tree_add_14_36_groupi_n_1854), .y(n_2504));
nand2 g53143 (.a(csa_tree_add_14_36_groupi_n_1854), .b(csa_tree_add_14_36_groupi_n_1834), .y(n_2506));
nand2 csa_tree_add_14_36_groupi_g53144 (.a(csa_tree_add_14_36_groupi_n_535), .b(csa_tree_add_14_36_groupi_n_350), .y(n_2507));
nand2 csa_tree_add_14_36_groupi_g53145 (.a(a_5), .b(b_15), .y(n_2508));
nand2 csa_tree_add_14_36_groupi_g53146 (.a(csa_tree_add_14_36_groupi_n_565), .b(csa_tree_add_14_36_groupi_n_428), .y(n_2509));
xor2 csa_tree_add_14_36_groupi_g51865__53147 (.a(n_2510), .b(n_2507), .y(n_2511));
xor2 csa_tree_add_14_36_groupi_g52120__53148 (.a(n_2509), .b(n_2508), .y(n_2510));
xor2 g67 (.a(n_2513), .b(csa_tree_add_14_36_groupi_n_741), .y(n_2514));
xor2 g68 (.a(n_2620), .b(csa_tree_add_14_36_groupi_n_101), .y(n_2513));
nand2 csa_tree_add_14_36_groupi_g53149 (.a(csa_tree_add_14_36_groupi_n_521), .b(csa_tree_add_14_36_groupi_n_354), .y(n_2515));
nand2 csa_tree_add_14_36_groupi_g53150 (.a(a_11), .b(b_15), .y(n_2516));
nand2 csa_tree_add_14_36_groupi_g53151 (.a(csa_tree_add_14_36_groupi_n_596), .b(csa_tree_add_14_36_groupi_n_449), .y(n_2517));
xor2 csa_tree_add_14_36_groupi_g51867__53152 (.a(n_2518), .b(n_2515), .y(n_2519));
xor2 csa_tree_add_14_36_groupi_g52117__53153 (.a(n_2517), .b(n_2516), .y(n_2518));
nand2 csa_tree_add_14_36_groupi_g53154 (.a(csa_tree_add_14_36_groupi_n_542), .b(csa_tree_add_14_36_groupi_n_319), .y(n_2520));
nand2 csa_tree_add_14_36_groupi_g53155 (.a(a_8), .b(b_15), .y(n_2521));
nand2 csa_tree_add_14_36_groupi_g53156 (.a(csa_tree_add_14_36_groupi_n_547), .b(csa_tree_add_14_36_groupi_n_427), .y(n_2522));
xor2 csa_tree_add_14_36_groupi_g51868__53157 (.a(n_2523), .b(n_2520), .y(n_2524));
xor2 csa_tree_add_14_36_groupi_g52119__53158 (.a(n_2522), .b(n_2521), .y(n_2523));
nand2 csa_tree_add_14_36_groupi_g53159 (.a(csa_tree_add_14_36_groupi_n_513), .b(csa_tree_add_14_36_groupi_n_409), .y(n_2525));
nand2 csa_tree_add_14_36_groupi_g53160 (.a(a_9), .b(b_15), .y(n_2526));
nand2 csa_tree_add_14_36_groupi_g53161 (.a(csa_tree_add_14_36_groupi_n_631), .b(csa_tree_add_14_36_groupi_n_450), .y(n_2527));
xor2 csa_tree_add_14_36_groupi_g51863__53162 (.a(n_2528), .b(n_2525), .y(n_2529));
xor2 csa_tree_add_14_36_groupi_g52121__53163 (.a(n_2527), .b(n_2526), .y(n_2528));
nor2 csa_tree_add_14_36_groupi_g53166 (.a(b_14), .b(b_13), .y(n_2537));
xor2 g57 (.a(n_2542), .b(csa_tree_add_14_36_groupi_n_1445), .y(n_2543));
xor2 g58 (.a(csa_tree_add_14_36_groupi_n_1338), .b(csa_tree_add_14_36_groupi_n_2064), .y(n_2542));
xor2 g59 (.a(csa_tree_add_14_36_groupi_n_1445), .b(csa_tree_add_14_36_groupi_n_1338), .y(n_2544));
nor2 g53168 (.a(n_2546), .b(n_2549), .y(n_2550));
inv g32 (.a(csa_tree_add_14_36_groupi_n_1651), .y(n_2546));
nand2 g28 (.a(csa_tree_add_14_36_groupi_n_1605), .b(n_2548), .y(n_2549));
inv g29 (.a(n_2547), .y(n_2548));
nand2 g30 (.a(csa_tree_add_14_36_groupi_n_2129), .b(csa_tree_add_14_36_groupi_n_2127), .y(n_2547));
nand2 g31 (.a(csa_tree_add_14_36_groupi_n_1651), .b(csa_tree_add_14_36_groupi_n_1605), .y(n_2551));
nand2 g53171 (.a(csa_tree_add_14_36_groupi_n_1013), .b(n_2553), .y(n_2554));
inv g53172 (.a(csa_tree_add_14_36_groupi_n_2108), .y(n_2553));
nand2 g53173 (.a(n_2634), .b(csa_tree_add_14_36_groupi_n_1013), .y(n_2556));
nand2 g53176 (.a(csa_tree_add_14_36_groupi_n_990), .b(n_2558), .y(n_2559));
inv g53177 (.a(csa_tree_add_14_36_groupi_n_2119), .y(n_2558));
nand2 g53178 (.a(n_2640), .b(csa_tree_add_14_36_groupi_n_990), .y(n_2561));
nand2 csa_tree_add_14_36_groupi_g51723__53179 (.a(csa_tree_add_14_36_groupi_n_1203), .b(csa_tree_add_14_36_groupi_n_1022), .y(n_2564));
xor2 csa_tree_add_14_36_groupi_g51568__53180 (.a(csa_tree_add_14_36_groupi_n_1285), .b(csa_tree_add_14_36_groupi_n_1216), .y(n_2565));
nand2 csa_tree_add_14_36_groupi_g51351__53181 (.a(n_2568), .b(csa_tree_add_14_36_groupi_n_1518), .y(n_2569));
xor2 csa_tree_add_14_36_groupi_g51432__53182 (.a(n_2567), .b(n_2564), .y(n_2568));
xor2 csa_tree_add_14_36_groupi_g51557__53183 (.a(n_2565), .b(n_2566), .y(n_2567));
inv csa_tree_add_14_36_groupi_g53184 (.a(csa_tree_add_14_36_groupi_n_1276), .y(n_2566));
nor2 csa_tree_add_14_36_groupi_g51350__53185 (.a(n_2568), .b(csa_tree_add_14_36_groupi_n_1518), .y(n_2570));
nor2 g53187 (.a(csa_tree_add_14_36_groupi_n_128), .b(n_2575), .y(n_2576));
nand2 g53189 (.a(b_9), .b(n_2574), .y(n_2575));
inv g53190 (.a(a_3), .y(n_2574));
nand2 g53191 (.a(csa_tree_add_14_36_groupi_n_129), .b(b_9), .y(n_2577));
nor2 g34 (.a(n_2582), .b(n_2585), .y(n_2586));
inv g38 (.a(csa_tree_add_14_36_groupi_n_465), .y(n_2582));
nand2 g35 (.a(csa_tree_add_14_36_groupi_n_99), .b(csa_tree_add_14_36_groupi_n_259), .y(n_2585));
inv g36 (.a(n_2583), .y(csa_tree_add_14_36_groupi_n_259));
xor2 g37 (.a(b_14), .b(b_13), .y(n_2583));
nand2 g53205 (.a(n_2606), .b(csa_tree_add_14_36_groupi_n_980), .y(n_2607));
inv g53206 (.a(n_2605), .y(n_2606));
xor2 g39 (.a(csa_tree_add_14_36_groupi_n_503), .b(csa_tree_add_14_36_groupi_n_2302), .y(n_2605));
nand2 g40 (.a(n_2645), .b(csa_tree_add_14_36_groupi_n_980), .y(n_2609));
nand2 g53209 (.a(csa_tree_add_14_36_groupi_n_979), .b(n_2611), .y(n_2612));
inv g53210 (.a(csa_tree_add_14_36_groupi_n_2128), .y(n_2611));
nand2 g53211 (.a(n_2657), .b(csa_tree_add_14_36_groupi_n_979), .y(n_2614));
nand2 g53212 (.a(b_14), .b(b_13), .y(n_2616));
nand2 g53213 (.a(n_2617), .b(b_9), .y(n_2618));
nand2 g53214 (.a(csa_tree_add_14_36_groupi_n_406), .b(csa_tree_add_14_36_groupi_n_255), .y(n_2617));
nand2 g11 (.a(n_2688), .b(b_3), .y(n_2620));
xor2 g71 (.a(csa_tree_add_14_36_groupi_n_1427), .b(n_2622), .y(n_2623));
xor2 g72 (.a(csa_tree_add_14_36_groupi_n_1189), .b(n_2621), .y(n_2622));
xor2 g73 (.a(csa_tree_add_14_36_groupi_n_1082), .b(csa_tree_add_14_36_groupi_n_1058), .y(n_2621));
xor2 g74 (.a(csa_tree_add_14_36_groupi_n_1427), .b(csa_tree_add_14_36_groupi_n_1189), .y(n_2624));
inv csa_tree_add_14_36_groupi_g53221 (.a(n_2633), .y(n_2634));
nor2 csa_tree_add_14_36_groupi_g51931__53222 (.a(n_2631), .b(n_2632), .y(n_2633));
nand2 csa_tree_add_14_36_groupi_g53223 (.a(n_157), .b(csa_tree_add_14_36_groupi_n_656), .y(n_2631));
nor2 csa_tree_add_14_36_groupi_g52029__53224 (.a(csa_tree_add_14_36_groupi_n_2116), .b(csa_tree_add_14_36_groupi_n_2054), .y(n_2632));
nor2 g53225 (.a(n_2633), .b(n_2554), .y(n_2635));
inv csa_tree_add_14_36_groupi_g53227 (.a(n_2639), .y(n_2640));
nor2 csa_tree_add_14_36_groupi_g51905__53228 (.a(n_2637), .b(n_2638), .y(n_2639));
nand2 csa_tree_add_14_36_groupi_g52165__53229 (.a(n_79), .b(csa_tree_add_14_36_groupi_n_2106), .y(n_2637));
nor2 csa_tree_add_14_36_groupi_g52021__53230 (.a(csa_tree_add_14_36_groupi_n_2073), .b(csa_tree_add_14_36_groupi_n_2062), .y(n_2638));
nor2 g53231 (.a(n_2639), .b(n_2559), .y(n_2641));
inv csa_tree_add_14_36_groupi_g53233 (.a(n_2644), .y(n_2645));
nor2 csa_tree_add_14_36_groupi_g51692__53234 (.a(n_2642), .b(n_2643), .y(n_2644));
nor2 csa_tree_add_14_36_groupi_g51884__53235 (.a(csa_tree_add_14_36_groupi_n_1071), .b(csa_tree_add_14_36_groupi_n_956), .y(n_2642));
nor2 csa_tree_add_14_36_groupi_g52062__53236 (.a(csa_tree_add_14_36_groupi_n_2140), .b(csa_tree_add_14_36_groupi_n_2092), .y(n_2643));
nor2 g53237 (.a(n_2644), .b(n_2607), .y(n_2646));
inv csa_tree_add_14_36_groupi_g53239 (.a(n_2656), .y(n_2657));
nor2 csa_tree_add_14_36_groupi_g51910__53240 (.a(n_2654), .b(n_2655), .y(n_2656));
nand2 csa_tree_add_14_36_groupi_g53241 (.a(n_77), .b(csa_tree_add_14_36_groupi_n_2123), .y(n_2654));
nor2 csa_tree_add_14_36_groupi_g52063__53242 (.a(csa_tree_add_14_36_groupi_n_2039), .b(csa_tree_add_14_36_groupi_n_2059), .y(n_2655));
nor2 g53243 (.a(n_2656), .b(n_2612), .y(n_2658));
xor2 g53245 (.a(b_11), .b(b_10), .y(n_2659));
inv g4 (.a(n_2674), .y(n_2675));
nor2 g53246 (.a(n_2673), .b(csa_tree_add_14_36_groupi_n_144), .y(n_2674));
nand2 csa_tree_add_14_36_groupi_g53247 (.a(n_2676), .b(n_2677), .y(n_2678));
inv csa_tree_add_14_36_groupi_g53248 (.a(csa_tree_add_14_36_groupi_n_144), .y(n_2676));
xor2 csa_tree_add_14_36_groupi_g53249 (.a(b_13), .b(b_12), .y(n_2677));
xor2 g53250 (.a(csa_tree_add_14_36_groupi_n_2254), .b(csa_tree_add_14_36_groupi_n_2219), .y(n_2681));
nand2 csa_tree_add_14_36_groupi_g51147__53251 (.a(n_2682), .b(csa_tree_add_14_36_groupi_n_2219), .y(n_2683));
inv csa_tree_add_14_36_groupi_g53252 (.a(csa_tree_add_14_36_groupi_n_2254), .y(n_2682));
nand2 csa_tree_add_14_36_groupi_g51142__53253 (.a(csa_tree_add_14_36_groupi_n_2254), .b(n_2684), .y(n_2685));
inv csa_tree_add_14_36_groupi_g53254 (.a(csa_tree_add_14_36_groupi_n_2219), .y(n_2684));
inv g53255 (.a(n_2687), .y(n_2688));
nor2 g53256 (.a(csa_tree_add_14_36_groupi_n_150), .b(csa_tree_add_14_36_groupi_n_230), .y(n_2687));
nand2 csa_tree_add_14_36_groupi_g53257 (.a(n_2689), .b(csa_tree_add_14_36_groupi_n_230), .y(n_2690));
inv csa_tree_add_14_36_groupi_g53258 (.a(csa_tree_add_14_36_groupi_n_150), .y(n_2689));
xor2 g53260 (.a(n_84), .b(csa_tree_add_14_36_groupi_n_2167), .y(n_2693));
nand2 csa_tree_add_14_36_groupi_g53261 (.a(n_2695), .b(csa_tree_add_14_36_groupi_n_2167), .y(n_2696));
inv csa_tree_add_14_36_groupi_g53262 (.a(n_84), .y(n_2695));
nand2 csa_tree_add_14_36_groupi_g53263 (.a(n_84), .b(n_2697), .y(n_2698));
inv csa_tree_add_14_36_groupi_g53264 (.a(csa_tree_add_14_36_groupi_n_2167), .y(n_2697));
inv g53282 (.a(b_12), .y(n_2673));
nor2 g304 (.a(n_2758), .b(n_2759), .y(n_2760));
nor2 g305 (.a(n_2756), .b(n_2757), .y(n_2758));
nand2 g306 (.a(n_2753), .b(n_2755), .y(n_2756));
nand2 g307 (.a(n_2751), .b(n_2752), .y(n_2753));
xor2 g310 (.a(n_2693), .b(csa_tree_add_14_36_groupi_n_2086), .y(n_2751));
nand2 g313 (.a(n_85), .b(csa_tree_add_14_36_groupi_n_2036), .y(n_2752));
inv g311 (.a(n_2754), .y(n_2755));
nor2 g312 (.a(csa_tree_add_14_36_groupi_n_498), .b(csa_tree_add_14_36_groupi_n_2135), .y(n_2754));
nor2 g314 (.a(csa_tree_add_14_36_groupi_n_891), .b(csa_tree_add_14_36_groupi_n_728), .y(n_2757));
nor2 g308 (.a(n_2751), .b(n_2752), .y(n_2759));
nor2 g309 (.a(n_2757), .b(n_2754), .y(n_2761));
nand2 g350 (.a(n_2769), .b(n_2770), .y(n_2771));
nand2 g351 (.a(n_2767), .b(n_2768), .y(n_2769));
inv g353 (.a(n_2766), .y(n_2767));
nor2 g354 (.a(n_2762), .b(n_2765), .y(n_2766));
xor2 g356 (.a(csa_tree_add_14_36_groupi_n_915), .b(csa_tree_add_14_36_groupi_n_725), .y(n_2762));
xor2 g355 (.a(n_2763), .b(n_2764), .y(n_2765));
xor2 g357 (.a(csa_tree_add_14_36_groupi_n_714), .b(csa_tree_add_14_36_groupi_n_718), .y(n_2763));
nand2 g359 (.a(csa_tree_add_14_36_groupi_n_634), .b(csa_tree_add_14_36_groupi_n_410), .y(n_2764));
nand2 g358 (.a(csa_tree_add_14_36_groupi_n_958), .b(csa_tree_add_14_36_groupi_n_861), .y(n_2768));
nand2 g352 (.a(n_2762), .b(n_2765), .y(n_2770));
nand2 g202 (.a(n_2774), .b(n_2777), .y(n_2778));
nand2 g205 (.a(n_2772), .b(csa_tree_add_14_36_groupi_n_80), .y(n_2774));
nand2 g207 (.a(n_151), .b(csa_tree_add_14_36_groupi_n_2043), .y(n_2772));
nor2 g204 (.a(n_2775), .b(n_2776), .y(n_2777));
nor2 g208 (.a(csa_tree_add_14_36_groupi_n_2102), .b(csa_tree_add_14_36_groupi_n_2094), .y(n_2775));
nor2 g210 (.a(n_151), .b(csa_tree_add_14_36_groupi_n_2043), .y(n_2776));
nand2 g203 (.a(n_2780), .b(n_2772), .y(n_2781));
nand2 g206 (.a(n_2779), .b(n_125), .y(n_2780));
inv g209 (.a(n_2776), .y(n_2779));
endmodule

